magic
tech sky130A
magscale 1 2
timestamp 1693011900
<< pwell >>
rect -352 -648 352 648
<< psubdiff >>
rect -316 578 -220 612
rect 220 578 316 612
rect -316 516 -282 578
rect 282 516 316 578
rect -316 -578 -282 -516
rect 282 -578 316 -516
rect -316 -612 -220 -578
rect 220 -612 316 -578
<< psubdiffcont >>
rect -220 578 220 612
rect -316 -516 -282 516
rect 282 -516 316 516
rect -220 -612 220 -578
<< xpolycontact >>
rect -186 50 -48 482
rect -186 -482 -48 -50
rect 48 50 186 482
rect 48 -482 186 -50
<< ppolyres >>
rect -186 -50 -48 50
rect 48 -50 186 50
<< locali >>
rect -316 578 -220 612
rect 220 578 316 612
rect -316 516 -282 578
rect 282 516 316 578
rect -316 -578 -282 -516
rect 282 -578 316 -516
rect -316 -612 -220 -578
rect 220 -612 316 -578
<< viali >>
rect -170 67 -64 464
rect 64 67 170 464
rect -170 -464 -64 -67
rect 64 -464 170 -67
<< metal1 >>
rect -176 464 -58 476
rect -176 67 -170 464
rect -64 67 -58 464
rect -176 55 -58 67
rect 58 464 176 476
rect 58 67 64 464
rect 170 67 176 464
rect 58 55 176 67
rect -176 -67 -58 -55
rect -176 -464 -170 -67
rect -64 -464 -58 -67
rect -176 -476 -58 -464
rect 58 -67 176 -55
rect 58 -464 64 -67
rect 170 -464 176 -67
rect 58 -476 176 -464
<< properties >>
string FIXED_BBOX -299 -595 299 595
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 0.50 m 1 nx 2 wmin 0.690 lmin 0.50 rho 319.8 val 796.434 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
