magic
tech sky130A
magscale 1 2
timestamp 1693420066
<< error_p >>
rect -1537 541 -1465 547
rect -1379 541 -1307 547
rect -1221 541 -1149 547
rect -1063 541 -991 547
rect -905 541 -833 547
rect -747 541 -675 547
rect -589 541 -517 547
rect -431 541 -359 547
rect -273 541 -201 547
rect -115 541 -43 547
rect 43 541 115 547
rect 201 541 273 547
rect 359 541 431 547
rect 517 541 589 547
rect 675 541 747 547
rect 833 541 905 547
rect 991 541 1063 547
rect 1149 541 1221 547
rect 1307 541 1379 547
rect 1465 541 1537 547
rect -1537 507 -1525 541
rect -1379 507 -1367 541
rect -1221 507 -1209 541
rect -1063 507 -1051 541
rect -905 507 -893 541
rect -747 507 -735 541
rect -589 507 -577 541
rect -431 507 -419 541
rect -273 507 -261 541
rect -115 507 -103 541
rect 43 507 55 541
rect 201 507 213 541
rect 359 507 371 541
rect 517 507 529 541
rect 675 507 687 541
rect 833 507 845 541
rect 991 507 1003 541
rect 1149 507 1161 541
rect 1307 507 1319 541
rect 1465 507 1477 541
rect -1537 501 -1465 507
rect -1379 501 -1307 507
rect -1221 501 -1149 507
rect -1063 501 -991 507
rect -905 501 -833 507
rect -747 501 -675 507
rect -589 501 -517 507
rect -431 501 -359 507
rect -273 501 -201 507
rect -115 501 -43 507
rect 43 501 115 507
rect 201 501 273 507
rect 359 501 431 507
rect 517 501 589 507
rect 675 501 747 507
rect 833 501 905 507
rect 991 501 1063 507
rect 1149 501 1221 507
rect 1307 501 1379 507
rect 1465 501 1537 507
<< pwell >>
rect -1779 -727 1779 727
<< mvnmos >>
rect -1551 -531 -1451 469
rect -1393 -531 -1293 469
rect -1235 -531 -1135 469
rect -1077 -531 -977 469
rect -919 -531 -819 469
rect -761 -531 -661 469
rect -603 -531 -503 469
rect -445 -531 -345 469
rect -287 -531 -187 469
rect -129 -531 -29 469
rect 29 -531 129 469
rect 187 -531 287 469
rect 345 -531 445 469
rect 503 -531 603 469
rect 661 -531 761 469
rect 819 -531 919 469
rect 977 -531 1077 469
rect 1135 -531 1235 469
rect 1293 -531 1393 469
rect 1451 -531 1551 469
<< mvndiff >>
rect -1609 457 -1551 469
rect -1609 -519 -1597 457
rect -1563 -519 -1551 457
rect -1609 -531 -1551 -519
rect -1451 457 -1393 469
rect -1451 -519 -1439 457
rect -1405 -519 -1393 457
rect -1451 -531 -1393 -519
rect -1293 457 -1235 469
rect -1293 -519 -1281 457
rect -1247 -519 -1235 457
rect -1293 -531 -1235 -519
rect -1135 457 -1077 469
rect -1135 -519 -1123 457
rect -1089 -519 -1077 457
rect -1135 -531 -1077 -519
rect -977 457 -919 469
rect -977 -519 -965 457
rect -931 -519 -919 457
rect -977 -531 -919 -519
rect -819 457 -761 469
rect -819 -519 -807 457
rect -773 -519 -761 457
rect -819 -531 -761 -519
rect -661 457 -603 469
rect -661 -519 -649 457
rect -615 -519 -603 457
rect -661 -531 -603 -519
rect -503 457 -445 469
rect -503 -519 -491 457
rect -457 -519 -445 457
rect -503 -531 -445 -519
rect -345 457 -287 469
rect -345 -519 -333 457
rect -299 -519 -287 457
rect -345 -531 -287 -519
rect -187 457 -129 469
rect -187 -519 -175 457
rect -141 -519 -129 457
rect -187 -531 -129 -519
rect -29 457 29 469
rect -29 -519 -17 457
rect 17 -519 29 457
rect -29 -531 29 -519
rect 129 457 187 469
rect 129 -519 141 457
rect 175 -519 187 457
rect 129 -531 187 -519
rect 287 457 345 469
rect 287 -519 299 457
rect 333 -519 345 457
rect 287 -531 345 -519
rect 445 457 503 469
rect 445 -519 457 457
rect 491 -519 503 457
rect 445 -531 503 -519
rect 603 457 661 469
rect 603 -519 615 457
rect 649 -519 661 457
rect 603 -531 661 -519
rect 761 457 819 469
rect 761 -519 773 457
rect 807 -519 819 457
rect 761 -531 819 -519
rect 919 457 977 469
rect 919 -519 931 457
rect 965 -519 977 457
rect 919 -531 977 -519
rect 1077 457 1135 469
rect 1077 -519 1089 457
rect 1123 -519 1135 457
rect 1077 -531 1135 -519
rect 1235 457 1293 469
rect 1235 -519 1247 457
rect 1281 -519 1293 457
rect 1235 -531 1293 -519
rect 1393 457 1451 469
rect 1393 -519 1405 457
rect 1439 -519 1451 457
rect 1393 -531 1451 -519
rect 1551 457 1609 469
rect 1551 -519 1563 457
rect 1597 -519 1609 457
rect 1551 -531 1609 -519
<< mvndiffc >>
rect -1597 -519 -1563 457
rect -1439 -519 -1405 457
rect -1281 -519 -1247 457
rect -1123 -519 -1089 457
rect -965 -519 -931 457
rect -807 -519 -773 457
rect -649 -519 -615 457
rect -491 -519 -457 457
rect -333 -519 -299 457
rect -175 -519 -141 457
rect -17 -519 17 457
rect 141 -519 175 457
rect 299 -519 333 457
rect 457 -519 491 457
rect 615 -519 649 457
rect 773 -519 807 457
rect 931 -519 965 457
rect 1089 -519 1123 457
rect 1247 -519 1281 457
rect 1405 -519 1439 457
rect 1563 -519 1597 457
<< mvpsubdiff >>
rect -1743 679 1743 691
rect -1743 645 -1635 679
rect 1635 645 1743 679
rect -1743 633 1743 645
rect -1743 583 -1685 633
rect -1743 -583 -1731 583
rect -1697 -583 -1685 583
rect 1685 583 1743 633
rect -1743 -633 -1685 -583
rect 1685 -583 1697 583
rect 1731 -583 1743 583
rect 1685 -633 1743 -583
rect -1743 -645 1743 -633
rect -1743 -679 -1635 -645
rect 1635 -679 1743 -645
rect -1743 -691 1743 -679
<< mvpsubdiffcont >>
rect -1635 645 1635 679
rect -1731 -583 -1697 583
rect 1697 -583 1731 583
rect -1635 -679 1635 -645
<< poly >>
rect -1537 541 -1465 557
rect -1537 524 -1521 541
rect -1551 507 -1521 524
rect -1481 524 -1465 541
rect -1379 541 -1307 557
rect -1379 524 -1363 541
rect -1481 507 -1451 524
rect -1551 469 -1451 507
rect -1393 507 -1363 524
rect -1323 524 -1307 541
rect -1221 541 -1149 557
rect -1221 524 -1205 541
rect -1323 507 -1293 524
rect -1393 469 -1293 507
rect -1235 507 -1205 524
rect -1165 524 -1149 541
rect -1063 541 -991 557
rect -1063 524 -1047 541
rect -1165 507 -1135 524
rect -1235 469 -1135 507
rect -1077 507 -1047 524
rect -1007 524 -991 541
rect -905 541 -833 557
rect -905 524 -889 541
rect -1007 507 -977 524
rect -1077 469 -977 507
rect -919 507 -889 524
rect -849 524 -833 541
rect -747 541 -675 557
rect -747 524 -731 541
rect -849 507 -819 524
rect -919 469 -819 507
rect -761 507 -731 524
rect -691 524 -675 541
rect -589 541 -517 557
rect -589 524 -573 541
rect -691 507 -661 524
rect -761 469 -661 507
rect -603 507 -573 524
rect -533 524 -517 541
rect -431 541 -359 557
rect -431 524 -415 541
rect -533 507 -503 524
rect -603 469 -503 507
rect -445 507 -415 524
rect -375 524 -359 541
rect -273 541 -201 557
rect -273 524 -257 541
rect -375 507 -345 524
rect -445 469 -345 507
rect -287 507 -257 524
rect -217 524 -201 541
rect -115 541 -43 557
rect -115 524 -99 541
rect -217 507 -187 524
rect -287 469 -187 507
rect -129 507 -99 524
rect -59 524 -43 541
rect 43 541 115 557
rect 43 524 59 541
rect -59 507 -29 524
rect -129 469 -29 507
rect 29 507 59 524
rect 99 524 115 541
rect 201 541 273 557
rect 201 524 217 541
rect 99 507 129 524
rect 29 469 129 507
rect 187 507 217 524
rect 257 524 273 541
rect 359 541 431 557
rect 359 524 375 541
rect 257 507 287 524
rect 187 469 287 507
rect 345 507 375 524
rect 415 524 431 541
rect 517 541 589 557
rect 517 524 533 541
rect 415 507 445 524
rect 345 469 445 507
rect 503 507 533 524
rect 573 524 589 541
rect 675 541 747 557
rect 675 524 691 541
rect 573 507 603 524
rect 503 469 603 507
rect 661 507 691 524
rect 731 524 747 541
rect 833 541 905 557
rect 833 524 849 541
rect 731 507 761 524
rect 661 469 761 507
rect 819 507 849 524
rect 889 524 905 541
rect 991 541 1063 557
rect 991 524 1007 541
rect 889 507 919 524
rect 819 469 919 507
rect 977 507 1007 524
rect 1047 524 1063 541
rect 1149 541 1221 557
rect 1149 524 1165 541
rect 1047 507 1077 524
rect 977 469 1077 507
rect 1135 507 1165 524
rect 1205 524 1221 541
rect 1307 541 1379 557
rect 1307 524 1323 541
rect 1205 507 1235 524
rect 1135 469 1235 507
rect 1293 507 1323 524
rect 1363 524 1379 541
rect 1465 541 1537 557
rect 1465 524 1481 541
rect 1363 507 1393 524
rect 1293 469 1393 507
rect 1451 507 1481 524
rect 1521 524 1537 541
rect 1521 507 1551 524
rect 1451 469 1551 507
rect -1551 -557 -1451 -531
rect -1393 -557 -1293 -531
rect -1235 -557 -1135 -531
rect -1077 -557 -977 -531
rect -919 -557 -819 -531
rect -761 -557 -661 -531
rect -603 -557 -503 -531
rect -445 -557 -345 -531
rect -287 -557 -187 -531
rect -129 -557 -29 -531
rect 29 -557 129 -531
rect 187 -557 287 -531
rect 345 -557 445 -531
rect 503 -557 603 -531
rect 661 -557 761 -531
rect 819 -557 919 -531
rect 977 -557 1077 -531
rect 1135 -557 1235 -531
rect 1293 -557 1393 -531
rect 1451 -557 1551 -531
<< polycont >>
rect -1521 507 -1481 541
rect -1363 507 -1323 541
rect -1205 507 -1165 541
rect -1047 507 -1007 541
rect -889 507 -849 541
rect -731 507 -691 541
rect -573 507 -533 541
rect -415 507 -375 541
rect -257 507 -217 541
rect -99 507 -59 541
rect 59 507 99 541
rect 217 507 257 541
rect 375 507 415 541
rect 533 507 573 541
rect 691 507 731 541
rect 849 507 889 541
rect 1007 507 1047 541
rect 1165 507 1205 541
rect 1323 507 1363 541
rect 1481 507 1521 541
<< locali >>
rect -1731 645 -1635 679
rect 1635 645 1731 679
rect -1731 583 -1697 645
rect 1697 583 1731 645
rect -1537 507 -1525 541
rect -1477 507 -1465 541
rect -1379 507 -1367 541
rect -1319 507 -1307 541
rect -1221 507 -1209 541
rect -1161 507 -1149 541
rect -1063 507 -1051 541
rect -1003 507 -991 541
rect -905 507 -893 541
rect -845 507 -833 541
rect -747 507 -735 541
rect -687 507 -675 541
rect -589 507 -577 541
rect -529 507 -517 541
rect -431 507 -419 541
rect -371 507 -359 541
rect -273 507 -261 541
rect -213 507 -201 541
rect -115 507 -103 541
rect -55 507 -43 541
rect 43 507 55 541
rect 103 507 115 541
rect 201 507 213 541
rect 261 507 273 541
rect 359 507 371 541
rect 419 507 431 541
rect 517 507 529 541
rect 577 507 589 541
rect 675 507 687 541
rect 735 507 747 541
rect 833 507 845 541
rect 893 507 905 541
rect 991 507 1003 541
rect 1051 507 1063 541
rect 1149 507 1161 541
rect 1209 507 1221 541
rect 1307 507 1319 541
rect 1367 507 1379 541
rect 1465 507 1477 541
rect 1525 507 1537 541
rect -1597 457 -1563 473
rect -1597 -535 -1563 -519
rect -1439 457 -1405 473
rect -1439 -535 -1405 -519
rect -1281 457 -1247 473
rect -1281 -535 -1247 -519
rect -1123 457 -1089 473
rect -1123 -535 -1089 -519
rect -965 457 -931 473
rect -965 -535 -931 -519
rect -807 457 -773 473
rect -807 -535 -773 -519
rect -649 457 -615 473
rect -649 -535 -615 -519
rect -491 457 -457 473
rect -491 -535 -457 -519
rect -333 457 -299 473
rect -333 -535 -299 -519
rect -175 457 -141 473
rect -175 -535 -141 -519
rect -17 457 17 473
rect -17 -535 17 -519
rect 141 457 175 473
rect 141 -535 175 -519
rect 299 457 333 473
rect 299 -535 333 -519
rect 457 457 491 473
rect 457 -535 491 -519
rect 615 457 649 473
rect 615 -535 649 -519
rect 773 457 807 473
rect 773 -535 807 -519
rect 931 457 965 473
rect 931 -535 965 -519
rect 1089 457 1123 473
rect 1089 -535 1123 -519
rect 1247 457 1281 473
rect 1247 -535 1281 -519
rect 1405 457 1439 473
rect 1405 -535 1439 -519
rect 1563 457 1597 473
rect 1563 -535 1597 -519
rect -1731 -645 -1697 -583
rect 1697 -645 1731 -583
rect -1731 -679 -1635 -645
rect 1635 -679 1731 -645
<< viali >>
rect -1525 507 -1521 541
rect -1521 507 -1481 541
rect -1481 507 -1477 541
rect -1367 507 -1363 541
rect -1363 507 -1323 541
rect -1323 507 -1319 541
rect -1209 507 -1205 541
rect -1205 507 -1165 541
rect -1165 507 -1161 541
rect -1051 507 -1047 541
rect -1047 507 -1007 541
rect -1007 507 -1003 541
rect -893 507 -889 541
rect -889 507 -849 541
rect -849 507 -845 541
rect -735 507 -731 541
rect -731 507 -691 541
rect -691 507 -687 541
rect -577 507 -573 541
rect -573 507 -533 541
rect -533 507 -529 541
rect -419 507 -415 541
rect -415 507 -375 541
rect -375 507 -371 541
rect -261 507 -257 541
rect -257 507 -217 541
rect -217 507 -213 541
rect -103 507 -99 541
rect -99 507 -59 541
rect -59 507 -55 541
rect 55 507 59 541
rect 59 507 99 541
rect 99 507 103 541
rect 213 507 217 541
rect 217 507 257 541
rect 257 507 261 541
rect 371 507 375 541
rect 375 507 415 541
rect 415 507 419 541
rect 529 507 533 541
rect 533 507 573 541
rect 573 507 577 541
rect 687 507 691 541
rect 691 507 731 541
rect 731 507 735 541
rect 845 507 849 541
rect 849 507 889 541
rect 889 507 893 541
rect 1003 507 1007 541
rect 1007 507 1047 541
rect 1047 507 1051 541
rect 1161 507 1165 541
rect 1165 507 1205 541
rect 1205 507 1209 541
rect 1319 507 1323 541
rect 1323 507 1363 541
rect 1363 507 1367 541
rect 1477 507 1481 541
rect 1481 507 1521 541
rect 1521 507 1525 541
rect -1597 -519 -1563 457
rect -1439 -519 -1405 457
rect -1281 -519 -1247 457
rect -1123 -519 -1089 457
rect -965 -519 -931 457
rect -807 -519 -773 457
rect -649 -519 -615 457
rect -491 -519 -457 457
rect -333 -519 -299 457
rect -175 -519 -141 457
rect -17 -519 17 457
rect 141 -519 175 457
rect 299 -519 333 457
rect 457 -519 491 457
rect 615 -519 649 457
rect 773 -519 807 457
rect 931 -519 965 457
rect 1089 -519 1123 457
rect 1247 -519 1281 457
rect 1405 -519 1439 457
rect 1563 -519 1597 457
<< metal1 >>
rect -1537 541 -1465 547
rect -1537 507 -1525 541
rect -1477 507 -1465 541
rect -1537 501 -1465 507
rect -1379 541 -1307 547
rect -1379 507 -1367 541
rect -1319 507 -1307 541
rect -1379 501 -1307 507
rect -1221 541 -1149 547
rect -1221 507 -1209 541
rect -1161 507 -1149 541
rect -1221 501 -1149 507
rect -1063 541 -991 547
rect -1063 507 -1051 541
rect -1003 507 -991 541
rect -1063 501 -991 507
rect -905 541 -833 547
rect -905 507 -893 541
rect -845 507 -833 541
rect -905 501 -833 507
rect -747 541 -675 547
rect -747 507 -735 541
rect -687 507 -675 541
rect -747 501 -675 507
rect -589 541 -517 547
rect -589 507 -577 541
rect -529 507 -517 541
rect -589 501 -517 507
rect -431 541 -359 547
rect -431 507 -419 541
rect -371 507 -359 541
rect -431 501 -359 507
rect -273 541 -201 547
rect -273 507 -261 541
rect -213 507 -201 541
rect -273 501 -201 507
rect -115 541 -43 547
rect -115 507 -103 541
rect -55 507 -43 541
rect -115 501 -43 507
rect 43 541 115 547
rect 43 507 55 541
rect 103 507 115 541
rect 43 501 115 507
rect 201 541 273 547
rect 201 507 213 541
rect 261 507 273 541
rect 201 501 273 507
rect 359 541 431 547
rect 359 507 371 541
rect 419 507 431 541
rect 359 501 431 507
rect 517 541 589 547
rect 517 507 529 541
rect 577 507 589 541
rect 517 501 589 507
rect 675 541 747 547
rect 675 507 687 541
rect 735 507 747 541
rect 675 501 747 507
rect 833 541 905 547
rect 833 507 845 541
rect 893 507 905 541
rect 833 501 905 507
rect 991 541 1063 547
rect 991 507 1003 541
rect 1051 507 1063 541
rect 991 501 1063 507
rect 1149 541 1221 547
rect 1149 507 1161 541
rect 1209 507 1221 541
rect 1149 501 1221 507
rect 1307 541 1379 547
rect 1307 507 1319 541
rect 1367 507 1379 541
rect 1307 501 1379 507
rect 1465 541 1537 547
rect 1465 507 1477 541
rect 1525 507 1537 541
rect 1465 501 1537 507
rect -1603 457 -1557 469
rect -1603 -519 -1597 457
rect -1563 -519 -1557 457
rect -1603 -531 -1557 -519
rect -1445 457 -1399 469
rect -1445 -519 -1439 457
rect -1405 -519 -1399 457
rect -1445 -531 -1399 -519
rect -1287 457 -1241 469
rect -1287 -519 -1281 457
rect -1247 -519 -1241 457
rect -1287 -531 -1241 -519
rect -1129 457 -1083 469
rect -1129 -519 -1123 457
rect -1089 -519 -1083 457
rect -1129 -531 -1083 -519
rect -971 457 -925 469
rect -971 -519 -965 457
rect -931 -519 -925 457
rect -971 -531 -925 -519
rect -813 457 -767 469
rect -813 -519 -807 457
rect -773 -519 -767 457
rect -813 -531 -767 -519
rect -655 457 -609 469
rect -655 -519 -649 457
rect -615 -519 -609 457
rect -655 -531 -609 -519
rect -497 457 -451 469
rect -497 -519 -491 457
rect -457 -519 -451 457
rect -497 -531 -451 -519
rect -339 457 -293 469
rect -339 -519 -333 457
rect -299 -519 -293 457
rect -339 -531 -293 -519
rect -181 457 -135 469
rect -181 -519 -175 457
rect -141 -519 -135 457
rect -181 -531 -135 -519
rect -23 457 23 469
rect -23 -519 -17 457
rect 17 -519 23 457
rect -23 -531 23 -519
rect 135 457 181 469
rect 135 -519 141 457
rect 175 -519 181 457
rect 135 -531 181 -519
rect 293 457 339 469
rect 293 -519 299 457
rect 333 -519 339 457
rect 293 -531 339 -519
rect 451 457 497 469
rect 451 -519 457 457
rect 491 -519 497 457
rect 451 -531 497 -519
rect 609 457 655 469
rect 609 -519 615 457
rect 649 -519 655 457
rect 609 -531 655 -519
rect 767 457 813 469
rect 767 -519 773 457
rect 807 -519 813 457
rect 767 -531 813 -519
rect 925 457 971 469
rect 925 -519 931 457
rect 965 -519 971 457
rect 925 -531 971 -519
rect 1083 457 1129 469
rect 1083 -519 1089 457
rect 1123 -519 1129 457
rect 1083 -531 1129 -519
rect 1241 457 1287 469
rect 1241 -519 1247 457
rect 1281 -519 1287 457
rect 1241 -531 1287 -519
rect 1399 457 1445 469
rect 1399 -519 1405 457
rect 1439 -519 1445 457
rect 1399 -531 1445 -519
rect 1557 457 1603 469
rect 1557 -519 1563 457
rect 1597 -519 1603 457
rect 1557 -531 1603 -519
<< properties >>
string FIXED_BBOX -1714 -662 1714 662
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.5 m 1 nf 20 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
