magic
tech sky130A
timestamp 1693418132
<< pwell >>
rect -443 -429 443 429
<< mvnmos >>
rect -329 -300 -129 300
rect -100 -300 100 300
rect 129 -300 329 300
<< mvndiff >>
rect -358 294 -329 300
rect -358 -294 -352 294
rect -335 -294 -329 294
rect -358 -300 -329 -294
rect -129 294 -100 300
rect -129 -294 -123 294
rect -106 -294 -100 294
rect -129 -300 -100 -294
rect 100 294 129 300
rect 100 -294 106 294
rect 123 -294 129 294
rect 100 -300 129 -294
rect 329 294 358 300
rect 329 -294 335 294
rect 352 -294 358 294
rect 329 -300 358 -294
<< mvndiffc >>
rect -352 -294 -335 294
rect -123 -294 -106 294
rect 106 -294 123 294
rect 335 -294 352 294
<< mvpsubdiff >>
rect -425 405 425 411
rect -425 388 -371 405
rect 371 388 425 405
rect -425 382 425 388
rect -425 357 -396 382
rect -425 -357 -419 357
rect -402 -357 -396 357
rect 396 357 425 382
rect -425 -382 -396 -357
rect 396 -357 402 357
rect 419 -357 425 357
rect 396 -382 425 -357
rect -425 -388 425 -382
rect -425 -405 -371 -388
rect 371 -405 425 -388
rect -425 -411 425 -405
<< mvpsubdiffcont >>
rect -371 388 371 405
rect -419 -357 -402 357
rect 402 -357 419 357
rect -371 -405 371 -388
<< poly >>
rect -329 336 -129 344
rect -329 319 -321 336
rect -137 319 -129 336
rect -329 300 -129 319
rect -100 336 100 344
rect -100 319 -92 336
rect 92 319 100 336
rect -100 300 100 319
rect 129 336 329 344
rect 129 319 137 336
rect 321 319 329 336
rect 129 300 329 319
rect -329 -319 -129 -300
rect -329 -336 -321 -319
rect -137 -336 -129 -319
rect -329 -344 -129 -336
rect -100 -319 100 -300
rect -100 -336 -92 -319
rect 92 -336 100 -319
rect -100 -344 100 -336
rect 129 -319 329 -300
rect 129 -336 137 -319
rect 321 -336 329 -319
rect 129 -344 329 -336
<< polycont >>
rect -321 319 -137 336
rect -92 319 92 336
rect 137 319 321 336
rect -321 -336 -137 -319
rect -92 -336 92 -319
rect 137 -336 321 -319
<< locali >>
rect -419 388 -371 405
rect 371 388 419 405
rect -419 357 -402 388
rect 402 357 419 388
rect -329 319 -321 336
rect -137 319 -129 336
rect -100 319 -92 336
rect 92 319 100 336
rect 129 319 137 336
rect 321 319 329 336
rect -352 294 -335 302
rect -352 -302 -335 -294
rect -123 294 -106 302
rect -123 -302 -106 -294
rect 106 294 123 302
rect 106 -302 123 -294
rect 335 294 352 302
rect 335 -302 352 -294
rect -329 -336 -321 -319
rect -137 -336 -129 -319
rect -100 -336 -92 -319
rect 92 -336 100 -319
rect 129 -336 137 -319
rect 321 -336 329 -319
rect -419 -388 -402 -357
rect 402 -388 419 -357
rect -419 -405 -371 -388
rect 371 -405 419 -388
<< viali >>
rect -321 319 -137 336
rect -92 319 92 336
rect 137 319 321 336
rect -352 -294 -335 294
rect -123 -294 -106 294
rect 106 -294 123 294
rect 335 -294 352 294
rect -321 -336 -137 -319
rect -92 -336 92 -319
rect 137 -336 321 -319
<< metal1 >>
rect -327 336 -131 339
rect -327 319 -321 336
rect -137 319 -131 336
rect -327 316 -131 319
rect -98 336 98 339
rect -98 319 -92 336
rect 92 319 98 336
rect -98 316 98 319
rect 131 336 327 339
rect 131 319 137 336
rect 321 319 327 336
rect 131 316 327 319
rect -355 294 -332 300
rect -355 -294 -352 294
rect -335 -294 -332 294
rect -355 -300 -332 -294
rect -126 294 -103 300
rect -126 -294 -123 294
rect -106 -294 -103 294
rect -126 -300 -103 -294
rect 103 294 126 300
rect 103 -294 106 294
rect 123 -294 126 294
rect 103 -300 126 -294
rect 332 294 355 300
rect 332 -294 335 294
rect 352 -294 355 294
rect 332 -300 355 -294
rect -327 -319 -131 -316
rect -327 -336 -321 -319
rect -137 -336 -131 -319
rect -327 -339 -131 -336
rect -98 -319 98 -316
rect -98 -336 -92 -319
rect 92 -336 98 -319
rect -98 -339 98 -336
rect 131 -319 327 -316
rect 131 -336 137 -319
rect 321 -336 327 -319
rect 131 -339 327 -336
<< properties >>
string FIXED_BBOX -410 -396 410 396
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 6 l 2 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
