* NGSPICE file created from cs_resistor_stage.ext - technology: sky130A

.subckt cs_resistor_stage_post VDD VSS VIN VOUT
X0 VSS VSS VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=0.87 ps=6.29 w=6 l=1
X1 VSS VIN VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X2 VSS VIN VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X3 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X4 VSS VIN VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X5 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X6 VSS VIN VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X7 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X8 VOUT VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.6 w=6 l=1
X9 VSS VIN VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X10 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X11 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X12 m1_682_1168# m1_516_78# VDD sky130_fd_pr__res_high_po_0p35 l=1
X13 VDD VDD VDD sky130_fd_pr__res_high_po_0p35 l=1
X14 m1_2176_1166# VOUT VDD sky130_fd_pr__res_high_po_0p35 l=1
X15 VDD VDD VDD sky130_fd_pr__res_high_po_0p35 l=1
X16 m1_848_1166# m1_1014_24# VDD sky130_fd_pr__res_high_po_0p35 l=1
X17 m1_2010_1168# m1_1844_78# VDD sky130_fd_pr__res_high_po_0p35 l=1
X18 VDD m1_516_78# VDD sky130_fd_pr__res_high_po_0p35 l=1
X19 m1_1346_1170# m1_1180_80# VDD sky130_fd_pr__res_high_po_0p35 l=1
X20 m1_1512_1166# m1_1014_24# VDD sky130_fd_pr__res_high_po_0p35 l=1
X21 m1_2010_1168# VOUT VDD sky130_fd_pr__res_high_po_0p35 l=1
X22 m1_1512_1166# m1_1678_22# VDD sky130_fd_pr__res_high_po_0p35 l=1
X23 m1_848_1166# m1_350_22# VDD sky130_fd_pr__res_high_po_0p35 l=1
X24 m1_682_1168# m1_1180_80# VDD sky130_fd_pr__res_high_po_0p35 l=1
X25 VDD m1_350_22# VDD sky130_fd_pr__res_high_po_0p35 l=1
X26 m1_2176_1166# m1_1678_22# VDD sky130_fd_pr__res_high_po_0p35 l=1
X27 m1_1346_1170# m1_1844_78# VDD sky130_fd_pr__res_high_po_0p35 l=1
C0 VIN m1_516_78# 0.00505f
C1 m1_2176_1166# VDD 0.121f
C2 m1_2010_1168# m1_1346_1170# 0.324f
C3 VIN VDD 0.287f
C4 m1_1512_1166# m1_848_1166# 1.94e-25
C5 m1_1014_24# m1_1512_1166# 0.0166f
C6 m1_1014_24# m1_848_1166# 0.0166f
C7 m1_350_22# m1_848_1166# 0.0166f
C8 m1_1678_22# m1_1512_1166# 0.0166f
C9 m1_2010_1168# VDD 0.513f
C10 m1_1014_24# m1_350_22# 0.324f
C11 VOUT VDD 0.646f
C12 m1_1014_24# m1_1678_22# 0.324f
C13 m1_1678_22# m1_350_22# 1.06e-19
C14 m1_1844_78# m1_1678_22# 0.744f
C15 m1_1180_80# m1_1346_1170# 0.0166f
C16 m1_1346_1170# m1_682_1168# 0.324f
C17 VIN m1_2176_1166# 0.00119f
C18 m1_516_78# m1_682_1168# 0.0166f
C19 m1_1180_80# VDD 0.12f
C20 m1_2010_1168# m1_2176_1166# 0.744f
C21 m1_682_1168# VDD 0.529f
C22 VOUT m1_2176_1166# 0.0201f
C23 VIN m1_2010_1168# 0.00112f
C24 VOUT VIN 3.23f
C25 m1_1346_1170# m1_1512_1166# 0.741f
C26 m1_1014_24# m1_1346_1170# 0.00423f
C27 VOUT m1_2010_1168# 0.0204f
C28 m1_1678_22# m1_1346_1170# 0.00423f
C29 m1_350_22# m1_516_78# 0.744f
C30 m1_1512_1166# VDD 0.121f
C31 VDD m1_848_1166# 0.121f
C32 m1_1844_78# m1_1346_1170# 0.0166f
C33 m1_1014_24# VDD 0.204f
C34 m1_350_22# VDD 0.534f
C35 m1_1678_22# VDD 0.205f
C36 m1_1844_78# VDD 0.121f
C37 VIN m1_1180_80# 0.00533f
C38 VIN m1_682_1168# 0.00128f
C39 VIN m1_1512_1166# 0.00108f
C40 VIN m1_848_1166# 0.0011f
C41 m1_1678_22# m1_2176_1166# 0.0166f
C42 m1_1014_24# VIN 0.00654f
C43 VIN m1_350_22# 0.008f
C44 m1_1678_22# VIN 0.008f
C45 VOUT m1_1512_1166# 0.00349f
C46 VOUT m1_848_1166# 0.00349f
C47 m1_1346_1170# VDD 0.206f
C48 m1_1014_24# VOUT 0.074f
C49 VOUT m1_350_22# 0.0744f
C50 m1_1844_78# VIN 0.00498f
C51 m1_1678_22# m1_2010_1168# 0.00423f
C52 m1_516_78# VDD 0.138f
C53 m1_1678_22# VOUT 0.399f
C54 m1_1180_80# m1_682_1168# 0.0166f
C55 m1_1844_78# m1_2010_1168# 0.0166f
C56 m1_682_1168# m1_848_1166# 0.744f
C57 m1_1014_24# m1_1180_80# 0.743f
C58 m1_1014_24# m1_682_1168# 0.00424f
C59 m1_350_22# m1_682_1168# 0.00423f
C60 VIN m1_1346_1170# 0.00128f
C61 m1_2176_1166# VSS 0.203f $ **FLOATING
C62 m1_2010_1168# VSS 0.314f $ **FLOATING
C63 m1_1844_78# VSS 0.207f $ **FLOATING
C64 m1_1678_22# VSS 0.236f $ **FLOATING
C65 m1_1512_1166# VSS 0.203f $ **FLOATING
C66 m1_1346_1170# VSS 0.303f $ **FLOATING
C67 m1_1180_80# VSS 0.207f $ **FLOATING
C68 m1_1014_24# VSS 0.236f $ **FLOATING
C69 m1_848_1166# VSS 0.203f $ **FLOATING
C70 m1_682_1168# VSS 0.303f $ **FLOATING
C71 m1_516_78# VSS 0.207f $ **FLOATING
C72 m1_350_22# VSS 0.246f $ **FLOATING
C73 VDD VSS 16.2f
C74 VOUT VSS 6.63f
C75 VIN VSS 6.19f
.ends
