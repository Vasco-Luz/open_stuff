magic
tech sky130A
magscale 1 2
timestamp 1693420540
<< locali >>
rect 116 126 152 740
rect 254 568 472 728
rect 2086 568 2304 710
rect 2406 126 2442 740
rect -20 -132 1438 20
rect 1582 -132 2578 20
rect -82 -300 -14 -132
rect 2920 -298 2990 -120
rect -144 -1462 -110 -1202
rect 3016 -1460 3050 -1200
<< viali >>
rect 1278 -1476 1470 -1442
<< metal1 >>
rect 1240 616 1320 800
rect 568 564 1846 616
rect 568 150 616 564
rect 1240 563 1320 564
rect 1026 100 1074 512
rect 1484 150 1532 564
rect 1942 100 1990 512
rect 1026 40 1990 100
rect 1438 -180 1582 40
rect 14 -210 2892 -180
rect -80 -300 -14 -236
rect 14 -242 48 -210
rect 84 -248 142 -242
rect 136 -300 142 -248
rect 84 -306 142 -300
rect 236 -248 300 -242
rect 236 -300 242 -248
rect 294 -300 300 -248
rect 236 -306 300 -300
rect 14 -358 48 -306
rect 330 -360 364 -210
rect 394 -248 458 -242
rect 394 -300 400 -248
rect 452 -300 458 -248
rect 394 -306 458 -300
rect 552 -248 616 -242
rect 552 -300 558 -248
rect 610 -300 616 -248
rect 552 -306 616 -300
rect 646 -358 680 -210
rect 710 -248 774 -242
rect 710 -300 716 -248
rect 768 -300 774 -248
rect 710 -306 774 -300
rect 868 -248 932 -242
rect 868 -300 874 -248
rect 926 -300 932 -248
rect 868 -306 932 -300
rect 962 -356 996 -210
rect 1026 -248 1090 -242
rect 1026 -300 1032 -248
rect 1084 -300 1090 -248
rect 1026 -306 1090 -300
rect 1184 -248 1248 -242
rect 1184 -300 1190 -248
rect 1242 -300 1248 -248
rect 1184 -306 1248 -300
rect 1278 -356 1312 -210
rect 1342 -248 1406 -242
rect 1342 -300 1348 -248
rect 1400 -300 1406 -248
rect 1342 -306 1406 -300
rect 1500 -248 1564 -242
rect 1500 -300 1506 -248
rect 1558 -300 1564 -248
rect 1500 -306 1564 -300
rect 1594 -358 1628 -210
rect 1658 -248 1722 -242
rect 1658 -300 1664 -248
rect 1716 -300 1722 -248
rect 1658 -306 1722 -300
rect 1816 -248 1880 -242
rect 1816 -300 1822 -248
rect 1874 -300 1880 -248
rect 1816 -306 1880 -300
rect 1910 -360 1944 -210
rect 1974 -248 2038 -242
rect 1974 -300 1980 -248
rect 2032 -300 2038 -248
rect 1974 -306 2038 -300
rect 2132 -248 2196 -242
rect 2132 -300 2138 -248
rect 2190 -300 2196 -248
rect 2132 -306 2196 -300
rect 2226 -354 2260 -210
rect 2290 -248 2354 -242
rect 2290 -300 2296 -248
rect 2348 -300 2354 -248
rect 2290 -306 2354 -300
rect 2448 -248 2512 -242
rect 2448 -300 2454 -248
rect 2506 -300 2512 -248
rect 2448 -306 2512 -300
rect 2542 -356 2576 -210
rect 2606 -248 2670 -242
rect 2606 -300 2612 -248
rect 2664 -300 2670 -248
rect 2606 -306 2670 -300
rect 2764 -248 2828 -242
rect 2764 -300 2770 -248
rect 2822 -300 2828 -248
rect 2764 -306 2828 -300
rect 2858 -358 2892 -210
rect 2920 -300 2988 -248
rect 172 -1380 206 -1326
rect 488 -1380 522 -1318
rect 804 -1380 838 -1316
rect 1120 -1380 1154 -1316
rect 1436 -1380 1470 -1314
rect 1752 -1380 1786 -1316
rect 2068 -1380 2102 -1318
rect 2384 -1380 2418 -1318
rect 2700 -1380 2734 -1318
rect 172 -1410 2734 -1380
rect 1266 -1442 1482 -1410
rect 1266 -1476 1278 -1442
rect 1470 -1476 1482 -1442
rect 1266 -1614 1482 -1476
<< via1 >>
rect 84 -300 136 -248
rect 242 -300 294 -248
rect 400 -300 452 -248
rect 558 -300 610 -248
rect 716 -300 768 -248
rect 874 -300 926 -248
rect 1032 -300 1084 -248
rect 1190 -300 1242 -248
rect 1348 -300 1400 -248
rect 1506 -300 1558 -248
rect 1664 -300 1716 -248
rect 1822 -300 1874 -248
rect 1980 -300 2032 -248
rect 2138 -300 2190 -248
rect 2296 -300 2348 -248
rect 2454 -300 2506 -248
rect 2612 -300 2664 -248
rect 2770 -300 2822 -248
<< metal2 >>
rect -378 -248 2828 -242
rect -378 -300 84 -248
rect 136 -300 242 -248
rect 294 -300 400 -248
rect 452 -300 558 -248
rect 610 -300 716 -248
rect 768 -300 874 -248
rect 926 -300 1032 -248
rect 1084 -300 1190 -248
rect 1242 -300 1348 -248
rect 1400 -300 1506 -248
rect 1558 -300 1664 -248
rect 1716 -300 1822 -248
rect 1874 -300 1980 -248
rect 2032 -300 2138 -248
rect 2190 -300 2296 -248
rect 2348 -300 2454 -248
rect 2506 -300 2612 -248
rect 2664 -300 2770 -248
rect 2822 -300 2828 -248
rect -378 -306 2828 -300
use sky130_fd_pr__nfet_g5v0d10v5_MQ566X  sky130_fd_pr__nfet_g5v0d10v5_MQ566X_0
timestamp 1693420066
transform 1 0 1453 0 1 -799
box -1779 -727 1779 727
use sky130_fd_pr__nfet_g5v0d10v5_QWVZXL  sky130_fd_pr__nfet_g5v0d10v5_QWVZXL_0
timestamp 1693418132
transform 1 0 1279 0 1 362
box -1344 -427 1344 427
<< labels >>
flabel metal1 1240 563 1320 800 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 1266 -1614 1482 -1476 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel metal2 -378 -306 84 -242 0 FreeSans 1600 0 0 0 VIN
port 5 nsew
flabel metal1 1438 -210 1582 100 0 FreeSans 1600 0 0 0 VOUT
port 7 nsew
<< end >>
