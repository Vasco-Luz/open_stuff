magic
tech sky130A
magscale 1 2
timestamp 1693012143
<< pwell >>
rect -1747 -6258 1747 6258
<< mvnmos >>
rect -1519 -6000 -1319 6000
rect -1261 -6000 -1061 6000
rect -1003 -6000 -803 6000
rect -745 -6000 -545 6000
rect -487 -6000 -287 6000
rect -229 -6000 -29 6000
rect 29 -6000 229 6000
rect 287 -6000 487 6000
rect 545 -6000 745 6000
rect 803 -6000 1003 6000
rect 1061 -6000 1261 6000
rect 1319 -6000 1519 6000
<< mvndiff >>
rect -1577 5988 -1519 6000
rect -1577 -5988 -1565 5988
rect -1531 -5988 -1519 5988
rect -1577 -6000 -1519 -5988
rect -1319 5988 -1261 6000
rect -1319 -5988 -1307 5988
rect -1273 -5988 -1261 5988
rect -1319 -6000 -1261 -5988
rect -1061 5988 -1003 6000
rect -1061 -5988 -1049 5988
rect -1015 -5988 -1003 5988
rect -1061 -6000 -1003 -5988
rect -803 5988 -745 6000
rect -803 -5988 -791 5988
rect -757 -5988 -745 5988
rect -803 -6000 -745 -5988
rect -545 5988 -487 6000
rect -545 -5988 -533 5988
rect -499 -5988 -487 5988
rect -545 -6000 -487 -5988
rect -287 5988 -229 6000
rect -287 -5988 -275 5988
rect -241 -5988 -229 5988
rect -287 -6000 -229 -5988
rect -29 5988 29 6000
rect -29 -5988 -17 5988
rect 17 -5988 29 5988
rect -29 -6000 29 -5988
rect 229 5988 287 6000
rect 229 -5988 241 5988
rect 275 -5988 287 5988
rect 229 -6000 287 -5988
rect 487 5988 545 6000
rect 487 -5988 499 5988
rect 533 -5988 545 5988
rect 487 -6000 545 -5988
rect 745 5988 803 6000
rect 745 -5988 757 5988
rect 791 -5988 803 5988
rect 745 -6000 803 -5988
rect 1003 5988 1061 6000
rect 1003 -5988 1015 5988
rect 1049 -5988 1061 5988
rect 1003 -6000 1061 -5988
rect 1261 5988 1319 6000
rect 1261 -5988 1273 5988
rect 1307 -5988 1319 5988
rect 1261 -6000 1319 -5988
rect 1519 5988 1577 6000
rect 1519 -5988 1531 5988
rect 1565 -5988 1577 5988
rect 1519 -6000 1577 -5988
<< mvndiffc >>
rect -1565 -5988 -1531 5988
rect -1307 -5988 -1273 5988
rect -1049 -5988 -1015 5988
rect -791 -5988 -757 5988
rect -533 -5988 -499 5988
rect -275 -5988 -241 5988
rect -17 -5988 17 5988
rect 241 -5988 275 5988
rect 499 -5988 533 5988
rect 757 -5988 791 5988
rect 1015 -5988 1049 5988
rect 1273 -5988 1307 5988
rect 1531 -5988 1565 5988
<< mvpsubdiff >>
rect -1711 6210 1711 6222
rect -1711 6176 -1603 6210
rect 1603 6176 1711 6210
rect -1711 6164 1711 6176
rect -1711 6114 -1653 6164
rect -1711 -6114 -1699 6114
rect -1665 -6114 -1653 6114
rect 1653 6114 1711 6164
rect -1711 -6164 -1653 -6114
rect 1653 -6114 1665 6114
rect 1699 -6114 1711 6114
rect 1653 -6164 1711 -6114
rect -1711 -6176 1711 -6164
rect -1711 -6210 -1603 -6176
rect 1603 -6210 1711 -6176
rect -1711 -6222 1711 -6210
<< mvpsubdiffcont >>
rect -1603 6176 1603 6210
rect -1699 -6114 -1665 6114
rect 1665 -6114 1699 6114
rect -1603 -6210 1603 -6176
<< poly >>
rect -1519 6072 -1319 6088
rect -1519 6038 -1503 6072
rect -1335 6038 -1319 6072
rect -1519 6000 -1319 6038
rect -1261 6072 -1061 6088
rect -1261 6038 -1245 6072
rect -1077 6038 -1061 6072
rect -1261 6000 -1061 6038
rect -1003 6072 -803 6088
rect -1003 6038 -987 6072
rect -819 6038 -803 6072
rect -1003 6000 -803 6038
rect -745 6072 -545 6088
rect -745 6038 -729 6072
rect -561 6038 -545 6072
rect -745 6000 -545 6038
rect -487 6072 -287 6088
rect -487 6038 -471 6072
rect -303 6038 -287 6072
rect -487 6000 -287 6038
rect -229 6072 -29 6088
rect -229 6038 -213 6072
rect -45 6038 -29 6072
rect -229 6000 -29 6038
rect 29 6072 229 6088
rect 29 6038 45 6072
rect 213 6038 229 6072
rect 29 6000 229 6038
rect 287 6072 487 6088
rect 287 6038 303 6072
rect 471 6038 487 6072
rect 287 6000 487 6038
rect 545 6072 745 6088
rect 545 6038 561 6072
rect 729 6038 745 6072
rect 545 6000 745 6038
rect 803 6072 1003 6088
rect 803 6038 819 6072
rect 987 6038 1003 6072
rect 803 6000 1003 6038
rect 1061 6072 1261 6088
rect 1061 6038 1077 6072
rect 1245 6038 1261 6072
rect 1061 6000 1261 6038
rect 1319 6072 1519 6088
rect 1319 6038 1335 6072
rect 1503 6038 1519 6072
rect 1319 6000 1519 6038
rect -1519 -6038 -1319 -6000
rect -1519 -6072 -1503 -6038
rect -1335 -6072 -1319 -6038
rect -1519 -6088 -1319 -6072
rect -1261 -6038 -1061 -6000
rect -1261 -6072 -1245 -6038
rect -1077 -6072 -1061 -6038
rect -1261 -6088 -1061 -6072
rect -1003 -6038 -803 -6000
rect -1003 -6072 -987 -6038
rect -819 -6072 -803 -6038
rect -1003 -6088 -803 -6072
rect -745 -6038 -545 -6000
rect -745 -6072 -729 -6038
rect -561 -6072 -545 -6038
rect -745 -6088 -545 -6072
rect -487 -6038 -287 -6000
rect -487 -6072 -471 -6038
rect -303 -6072 -287 -6038
rect -487 -6088 -287 -6072
rect -229 -6038 -29 -6000
rect -229 -6072 -213 -6038
rect -45 -6072 -29 -6038
rect -229 -6088 -29 -6072
rect 29 -6038 229 -6000
rect 29 -6072 45 -6038
rect 213 -6072 229 -6038
rect 29 -6088 229 -6072
rect 287 -6038 487 -6000
rect 287 -6072 303 -6038
rect 471 -6072 487 -6038
rect 287 -6088 487 -6072
rect 545 -6038 745 -6000
rect 545 -6072 561 -6038
rect 729 -6072 745 -6038
rect 545 -6088 745 -6072
rect 803 -6038 1003 -6000
rect 803 -6072 819 -6038
rect 987 -6072 1003 -6038
rect 803 -6088 1003 -6072
rect 1061 -6038 1261 -6000
rect 1061 -6072 1077 -6038
rect 1245 -6072 1261 -6038
rect 1061 -6088 1261 -6072
rect 1319 -6038 1519 -6000
rect 1319 -6072 1335 -6038
rect 1503 -6072 1519 -6038
rect 1319 -6088 1519 -6072
<< polycont >>
rect -1503 6038 -1335 6072
rect -1245 6038 -1077 6072
rect -987 6038 -819 6072
rect -729 6038 -561 6072
rect -471 6038 -303 6072
rect -213 6038 -45 6072
rect 45 6038 213 6072
rect 303 6038 471 6072
rect 561 6038 729 6072
rect 819 6038 987 6072
rect 1077 6038 1245 6072
rect 1335 6038 1503 6072
rect -1503 -6072 -1335 -6038
rect -1245 -6072 -1077 -6038
rect -987 -6072 -819 -6038
rect -729 -6072 -561 -6038
rect -471 -6072 -303 -6038
rect -213 -6072 -45 -6038
rect 45 -6072 213 -6038
rect 303 -6072 471 -6038
rect 561 -6072 729 -6038
rect 819 -6072 987 -6038
rect 1077 -6072 1245 -6038
rect 1335 -6072 1503 -6038
<< locali >>
rect -1699 6176 -1603 6210
rect 1603 6176 1699 6210
rect -1699 6114 -1665 6176
rect 1665 6114 1699 6176
rect -1519 6038 -1503 6072
rect -1335 6038 -1319 6072
rect -1261 6038 -1245 6072
rect -1077 6038 -1061 6072
rect -1003 6038 -987 6072
rect -819 6038 -803 6072
rect -745 6038 -729 6072
rect -561 6038 -545 6072
rect -487 6038 -471 6072
rect -303 6038 -287 6072
rect -229 6038 -213 6072
rect -45 6038 -29 6072
rect 29 6038 45 6072
rect 213 6038 229 6072
rect 287 6038 303 6072
rect 471 6038 487 6072
rect 545 6038 561 6072
rect 729 6038 745 6072
rect 803 6038 819 6072
rect 987 6038 1003 6072
rect 1061 6038 1077 6072
rect 1245 6038 1261 6072
rect 1319 6038 1335 6072
rect 1503 6038 1519 6072
rect -1565 5988 -1531 6004
rect -1565 -6004 -1531 -5988
rect -1307 5988 -1273 6004
rect -1307 -6004 -1273 -5988
rect -1049 5988 -1015 6004
rect -1049 -6004 -1015 -5988
rect -791 5988 -757 6004
rect -791 -6004 -757 -5988
rect -533 5988 -499 6004
rect -533 -6004 -499 -5988
rect -275 5988 -241 6004
rect -275 -6004 -241 -5988
rect -17 5988 17 6004
rect -17 -6004 17 -5988
rect 241 5988 275 6004
rect 241 -6004 275 -5988
rect 499 5988 533 6004
rect 499 -6004 533 -5988
rect 757 5988 791 6004
rect 757 -6004 791 -5988
rect 1015 5988 1049 6004
rect 1015 -6004 1049 -5988
rect 1273 5988 1307 6004
rect 1273 -6004 1307 -5988
rect 1531 5988 1565 6004
rect 1531 -6004 1565 -5988
rect -1519 -6072 -1503 -6038
rect -1335 -6072 -1319 -6038
rect -1261 -6072 -1245 -6038
rect -1077 -6072 -1061 -6038
rect -1003 -6072 -987 -6038
rect -819 -6072 -803 -6038
rect -745 -6072 -729 -6038
rect -561 -6072 -545 -6038
rect -487 -6072 -471 -6038
rect -303 -6072 -287 -6038
rect -229 -6072 -213 -6038
rect -45 -6072 -29 -6038
rect 29 -6072 45 -6038
rect 213 -6072 229 -6038
rect 287 -6072 303 -6038
rect 471 -6072 487 -6038
rect 545 -6072 561 -6038
rect 729 -6072 745 -6038
rect 803 -6072 819 -6038
rect 987 -6072 1003 -6038
rect 1061 -6072 1077 -6038
rect 1245 -6072 1261 -6038
rect 1319 -6072 1335 -6038
rect 1503 -6072 1519 -6038
rect -1699 -6176 -1665 -6114
rect 1665 -6176 1699 -6114
rect -1699 -6210 -1603 -6176
rect 1603 -6210 1699 -6176
<< viali >>
rect -1503 6038 -1335 6072
rect -1245 6038 -1077 6072
rect -987 6038 -819 6072
rect -729 6038 -561 6072
rect -471 6038 -303 6072
rect -213 6038 -45 6072
rect 45 6038 213 6072
rect 303 6038 471 6072
rect 561 6038 729 6072
rect 819 6038 987 6072
rect 1077 6038 1245 6072
rect 1335 6038 1503 6072
rect -1565 -5988 -1531 5988
rect -1307 -5988 -1273 5988
rect -1049 -5988 -1015 5988
rect -791 -5988 -757 5988
rect -533 -5988 -499 5988
rect -275 -5988 -241 5988
rect -17 -5988 17 5988
rect 241 -5988 275 5988
rect 499 -5988 533 5988
rect 757 -5988 791 5988
rect 1015 -5988 1049 5988
rect 1273 -5988 1307 5988
rect 1531 -5988 1565 5988
rect -1503 -6072 -1335 -6038
rect -1245 -6072 -1077 -6038
rect -987 -6072 -819 -6038
rect -729 -6072 -561 -6038
rect -471 -6072 -303 -6038
rect -213 -6072 -45 -6038
rect 45 -6072 213 -6038
rect 303 -6072 471 -6038
rect 561 -6072 729 -6038
rect 819 -6072 987 -6038
rect 1077 -6072 1245 -6038
rect 1335 -6072 1503 -6038
<< metal1 >>
rect -1515 6072 -1323 6078
rect -1515 6038 -1503 6072
rect -1335 6038 -1323 6072
rect -1515 6032 -1323 6038
rect -1257 6072 -1065 6078
rect -1257 6038 -1245 6072
rect -1077 6038 -1065 6072
rect -1257 6032 -1065 6038
rect -999 6072 -807 6078
rect -999 6038 -987 6072
rect -819 6038 -807 6072
rect -999 6032 -807 6038
rect -741 6072 -549 6078
rect -741 6038 -729 6072
rect -561 6038 -549 6072
rect -741 6032 -549 6038
rect -483 6072 -291 6078
rect -483 6038 -471 6072
rect -303 6038 -291 6072
rect -483 6032 -291 6038
rect -225 6072 -33 6078
rect -225 6038 -213 6072
rect -45 6038 -33 6072
rect -225 6032 -33 6038
rect 33 6072 225 6078
rect 33 6038 45 6072
rect 213 6038 225 6072
rect 33 6032 225 6038
rect 291 6072 483 6078
rect 291 6038 303 6072
rect 471 6038 483 6072
rect 291 6032 483 6038
rect 549 6072 741 6078
rect 549 6038 561 6072
rect 729 6038 741 6072
rect 549 6032 741 6038
rect 807 6072 999 6078
rect 807 6038 819 6072
rect 987 6038 999 6072
rect 807 6032 999 6038
rect 1065 6072 1257 6078
rect 1065 6038 1077 6072
rect 1245 6038 1257 6072
rect 1065 6032 1257 6038
rect 1323 6072 1515 6078
rect 1323 6038 1335 6072
rect 1503 6038 1515 6072
rect 1323 6032 1515 6038
rect -1571 5988 -1525 6000
rect -1571 -5988 -1565 5988
rect -1531 -5988 -1525 5988
rect -1571 -6000 -1525 -5988
rect -1313 5988 -1267 6000
rect -1313 -5988 -1307 5988
rect -1273 -5988 -1267 5988
rect -1313 -6000 -1267 -5988
rect -1055 5988 -1009 6000
rect -1055 -5988 -1049 5988
rect -1015 -5988 -1009 5988
rect -1055 -6000 -1009 -5988
rect -797 5988 -751 6000
rect -797 -5988 -791 5988
rect -757 -5988 -751 5988
rect -797 -6000 -751 -5988
rect -539 5988 -493 6000
rect -539 -5988 -533 5988
rect -499 -5988 -493 5988
rect -539 -6000 -493 -5988
rect -281 5988 -235 6000
rect -281 -5988 -275 5988
rect -241 -5988 -235 5988
rect -281 -6000 -235 -5988
rect -23 5988 23 6000
rect -23 -5988 -17 5988
rect 17 -5988 23 5988
rect -23 -6000 23 -5988
rect 235 5988 281 6000
rect 235 -5988 241 5988
rect 275 -5988 281 5988
rect 235 -6000 281 -5988
rect 493 5988 539 6000
rect 493 -5988 499 5988
rect 533 -5988 539 5988
rect 493 -6000 539 -5988
rect 751 5988 797 6000
rect 751 -5988 757 5988
rect 791 -5988 797 5988
rect 751 -6000 797 -5988
rect 1009 5988 1055 6000
rect 1009 -5988 1015 5988
rect 1049 -5988 1055 5988
rect 1009 -6000 1055 -5988
rect 1267 5988 1313 6000
rect 1267 -5988 1273 5988
rect 1307 -5988 1313 5988
rect 1267 -6000 1313 -5988
rect 1525 5988 1571 6000
rect 1525 -5988 1531 5988
rect 1565 -5988 1571 5988
rect 1525 -6000 1571 -5988
rect -1515 -6038 -1323 -6032
rect -1515 -6072 -1503 -6038
rect -1335 -6072 -1323 -6038
rect -1515 -6078 -1323 -6072
rect -1257 -6038 -1065 -6032
rect -1257 -6072 -1245 -6038
rect -1077 -6072 -1065 -6038
rect -1257 -6078 -1065 -6072
rect -999 -6038 -807 -6032
rect -999 -6072 -987 -6038
rect -819 -6072 -807 -6038
rect -999 -6078 -807 -6072
rect -741 -6038 -549 -6032
rect -741 -6072 -729 -6038
rect -561 -6072 -549 -6038
rect -741 -6078 -549 -6072
rect -483 -6038 -291 -6032
rect -483 -6072 -471 -6038
rect -303 -6072 -291 -6038
rect -483 -6078 -291 -6072
rect -225 -6038 -33 -6032
rect -225 -6072 -213 -6038
rect -45 -6072 -33 -6038
rect -225 -6078 -33 -6072
rect 33 -6038 225 -6032
rect 33 -6072 45 -6038
rect 213 -6072 225 -6038
rect 33 -6078 225 -6072
rect 291 -6038 483 -6032
rect 291 -6072 303 -6038
rect 471 -6072 483 -6038
rect 291 -6078 483 -6072
rect 549 -6038 741 -6032
rect 549 -6072 561 -6038
rect 729 -6072 741 -6038
rect 549 -6078 741 -6072
rect 807 -6038 999 -6032
rect 807 -6072 819 -6038
rect 987 -6072 999 -6038
rect 807 -6078 999 -6072
rect 1065 -6038 1257 -6032
rect 1065 -6072 1077 -6038
rect 1245 -6072 1257 -6038
rect 1065 -6078 1257 -6072
rect 1323 -6038 1515 -6032
rect 1323 -6072 1335 -6038
rect 1503 -6072 1515 -6038
rect 1323 -6078 1515 -6072
<< properties >>
string FIXED_BBOX -1682 -6193 1682 6193
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 60 l 1 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
