magic
tech sky130A
magscale 1 2
timestamp 1693264311
<< pwell >>
rect -1612 -698 1612 698
<< psubdiff >>
rect -1576 628 -1480 662
rect 1480 628 1576 662
rect -1576 566 -1542 628
rect 1542 566 1576 628
rect -1576 -628 -1542 -566
rect 1542 -628 1576 -566
rect -1576 -662 -1480 -628
rect 1480 -662 1576 -628
<< psubdiffcont >>
rect -1480 628 1480 662
rect -1576 -566 -1542 566
rect 1542 -566 1576 566
rect -1480 -662 1480 -628
<< xpolycontact >>
rect -1446 100 -1376 532
rect -1446 -532 -1376 -100
rect -1280 100 -1210 532
rect -1280 -532 -1210 -100
rect -1114 100 -1044 532
rect -1114 -532 -1044 -100
rect -948 100 -878 532
rect -948 -532 -878 -100
rect -782 100 -712 532
rect -782 -532 -712 -100
rect -616 100 -546 532
rect -616 -532 -546 -100
rect -450 100 -380 532
rect -450 -532 -380 -100
rect -284 100 -214 532
rect -284 -532 -214 -100
rect -118 100 -48 532
rect -118 -532 -48 -100
rect 48 100 118 532
rect 48 -532 118 -100
rect 214 100 284 532
rect 214 -532 284 -100
rect 380 100 450 532
rect 380 -532 450 -100
rect 546 100 616 532
rect 546 -532 616 -100
rect 712 100 782 532
rect 712 -532 782 -100
rect 878 100 948 532
rect 878 -532 948 -100
rect 1044 100 1114 532
rect 1044 -532 1114 -100
rect 1210 100 1280 532
rect 1210 -532 1280 -100
rect 1376 100 1446 532
rect 1376 -532 1446 -100
<< ppolyres >>
rect -1446 -100 -1376 100
rect -1280 -100 -1210 100
rect -1114 -100 -1044 100
rect -948 -100 -878 100
rect -782 -100 -712 100
rect -616 -100 -546 100
rect -450 -100 -380 100
rect -284 -100 -214 100
rect -118 -100 -48 100
rect 48 -100 118 100
rect 214 -100 284 100
rect 380 -100 450 100
rect 546 -100 616 100
rect 712 -100 782 100
rect 878 -100 948 100
rect 1044 -100 1114 100
rect 1210 -100 1280 100
rect 1376 -100 1446 100
<< locali >>
rect -1576 628 -1480 662
rect 1480 628 1576 662
rect -1576 566 -1542 628
rect 1542 566 1576 628
rect -1576 -628 -1542 -566
rect 1542 -628 1576 -566
rect -1576 -662 -1480 -628
rect 1480 -662 1576 -628
<< viali >>
rect -1430 117 -1392 514
rect -1264 117 -1226 514
rect -1098 117 -1060 514
rect -932 117 -894 514
rect -766 117 -728 514
rect -600 117 -562 514
rect -434 117 -396 514
rect -268 117 -230 514
rect -102 117 -64 514
rect 64 117 102 514
rect 230 117 268 514
rect 396 117 434 514
rect 562 117 600 514
rect 728 117 766 514
rect 894 117 932 514
rect 1060 117 1098 514
rect 1226 117 1264 514
rect 1392 117 1430 514
rect -1430 -514 -1392 -117
rect -1264 -514 -1226 -117
rect -1098 -514 -1060 -117
rect -932 -514 -894 -117
rect -766 -514 -728 -117
rect -600 -514 -562 -117
rect -434 -514 -396 -117
rect -268 -514 -230 -117
rect -102 -514 -64 -117
rect 64 -514 102 -117
rect 230 -514 268 -117
rect 396 -514 434 -117
rect 562 -514 600 -117
rect 728 -514 766 -117
rect 894 -514 932 -117
rect 1060 -514 1098 -117
rect 1226 -514 1264 -117
rect 1392 -514 1430 -117
<< metal1 >>
rect -1436 514 -1386 526
rect -1436 117 -1430 514
rect -1392 117 -1386 514
rect -1436 105 -1386 117
rect -1270 514 -1220 526
rect -1270 117 -1264 514
rect -1226 117 -1220 514
rect -1270 105 -1220 117
rect -1104 514 -1054 526
rect -1104 117 -1098 514
rect -1060 117 -1054 514
rect -1104 105 -1054 117
rect -938 514 -888 526
rect -938 117 -932 514
rect -894 117 -888 514
rect -938 105 -888 117
rect -772 514 -722 526
rect -772 117 -766 514
rect -728 117 -722 514
rect -772 105 -722 117
rect -606 514 -556 526
rect -606 117 -600 514
rect -562 117 -556 514
rect -606 105 -556 117
rect -440 514 -390 526
rect -440 117 -434 514
rect -396 117 -390 514
rect -440 105 -390 117
rect -274 514 -224 526
rect -274 117 -268 514
rect -230 117 -224 514
rect -274 105 -224 117
rect -108 514 -58 526
rect -108 117 -102 514
rect -64 117 -58 514
rect -108 105 -58 117
rect 58 514 108 526
rect 58 117 64 514
rect 102 117 108 514
rect 58 105 108 117
rect 224 514 274 526
rect 224 117 230 514
rect 268 117 274 514
rect 224 105 274 117
rect 390 514 440 526
rect 390 117 396 514
rect 434 117 440 514
rect 390 105 440 117
rect 556 514 606 526
rect 556 117 562 514
rect 600 117 606 514
rect 556 105 606 117
rect 722 514 772 526
rect 722 117 728 514
rect 766 117 772 514
rect 722 105 772 117
rect 888 514 938 526
rect 888 117 894 514
rect 932 117 938 514
rect 888 105 938 117
rect 1054 514 1104 526
rect 1054 117 1060 514
rect 1098 117 1104 514
rect 1054 105 1104 117
rect 1220 514 1270 526
rect 1220 117 1226 514
rect 1264 117 1270 514
rect 1220 105 1270 117
rect 1386 514 1436 526
rect 1386 117 1392 514
rect 1430 117 1436 514
rect 1386 105 1436 117
rect -1436 -117 -1386 -105
rect -1436 -514 -1430 -117
rect -1392 -514 -1386 -117
rect -1436 -526 -1386 -514
rect -1270 -117 -1220 -105
rect -1270 -514 -1264 -117
rect -1226 -514 -1220 -117
rect -1270 -526 -1220 -514
rect -1104 -117 -1054 -105
rect -1104 -514 -1098 -117
rect -1060 -514 -1054 -117
rect -1104 -526 -1054 -514
rect -938 -117 -888 -105
rect -938 -514 -932 -117
rect -894 -514 -888 -117
rect -938 -526 -888 -514
rect -772 -117 -722 -105
rect -772 -514 -766 -117
rect -728 -514 -722 -117
rect -772 -526 -722 -514
rect -606 -117 -556 -105
rect -606 -514 -600 -117
rect -562 -514 -556 -117
rect -606 -526 -556 -514
rect -440 -117 -390 -105
rect -440 -514 -434 -117
rect -396 -514 -390 -117
rect -440 -526 -390 -514
rect -274 -117 -224 -105
rect -274 -514 -268 -117
rect -230 -514 -224 -117
rect -274 -526 -224 -514
rect -108 -117 -58 -105
rect -108 -514 -102 -117
rect -64 -514 -58 -117
rect -108 -526 -58 -514
rect 58 -117 108 -105
rect 58 -514 64 -117
rect 102 -514 108 -117
rect 58 -526 108 -514
rect 224 -117 274 -105
rect 224 -514 230 -117
rect 268 -514 274 -117
rect 224 -526 274 -514
rect 390 -117 440 -105
rect 390 -514 396 -117
rect 434 -514 440 -117
rect 390 -526 440 -514
rect 556 -117 606 -105
rect 556 -514 562 -117
rect 600 -514 606 -117
rect 556 -526 606 -514
rect 722 -117 772 -105
rect 722 -514 728 -117
rect 766 -514 772 -117
rect 722 -526 772 -514
rect 888 -117 938 -105
rect 888 -514 894 -117
rect 932 -514 938 -117
rect 888 -526 938 -514
rect 1054 -117 1104 -105
rect 1054 -514 1060 -117
rect 1098 -514 1104 -117
rect 1054 -526 1104 -514
rect 1220 -117 1270 -105
rect 1220 -514 1226 -117
rect 1264 -514 1270 -117
rect 1220 -526 1270 -514
rect 1386 -117 1436 -105
rect 1386 -514 1392 -117
rect 1430 -514 1436 -117
rect 1386 -526 1436 -514
<< properties >>
string FIXED_BBOX -1559 -645 1559 645
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.35 l 1.0 m 1 nx 18 wmin 0.350 lmin 0.50 rho 319.8 val 2.026k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
