magic
tech sky130A
magscale 1 2
timestamp 1693046372
<< pwell >>
rect -1747 -827 1747 827
<< mvnmos >>
rect -1519 -631 -1319 569
rect -1261 -631 -1061 569
rect -1003 -631 -803 569
rect -745 -631 -545 569
rect -487 -631 -287 569
rect -229 -631 -29 569
rect 29 -631 229 569
rect 287 -631 487 569
rect 545 -631 745 569
rect 803 -631 1003 569
rect 1061 -631 1261 569
rect 1319 -631 1519 569
<< mvndiff >>
rect -1577 557 -1519 569
rect -1577 -619 -1565 557
rect -1531 -619 -1519 557
rect -1577 -631 -1519 -619
rect -1319 557 -1261 569
rect -1319 -619 -1307 557
rect -1273 -619 -1261 557
rect -1319 -631 -1261 -619
rect -1061 557 -1003 569
rect -1061 -619 -1049 557
rect -1015 -619 -1003 557
rect -1061 -631 -1003 -619
rect -803 557 -745 569
rect -803 -619 -791 557
rect -757 -619 -745 557
rect -803 -631 -745 -619
rect -545 557 -487 569
rect -545 -619 -533 557
rect -499 -619 -487 557
rect -545 -631 -487 -619
rect -287 557 -229 569
rect -287 -619 -275 557
rect -241 -619 -229 557
rect -287 -631 -229 -619
rect -29 557 29 569
rect -29 -619 -17 557
rect 17 -619 29 557
rect -29 -631 29 -619
rect 229 557 287 569
rect 229 -619 241 557
rect 275 -619 287 557
rect 229 -631 287 -619
rect 487 557 545 569
rect 487 -619 499 557
rect 533 -619 545 557
rect 487 -631 545 -619
rect 745 557 803 569
rect 745 -619 757 557
rect 791 -619 803 557
rect 745 -631 803 -619
rect 1003 557 1061 569
rect 1003 -619 1015 557
rect 1049 -619 1061 557
rect 1003 -631 1061 -619
rect 1261 557 1319 569
rect 1261 -619 1273 557
rect 1307 -619 1319 557
rect 1261 -631 1319 -619
rect 1519 557 1577 569
rect 1519 -619 1531 557
rect 1565 -619 1577 557
rect 1519 -631 1577 -619
<< mvndiffc >>
rect -1565 -619 -1531 557
rect -1307 -619 -1273 557
rect -1049 -619 -1015 557
rect -791 -619 -757 557
rect -533 -619 -499 557
rect -275 -619 -241 557
rect -17 -619 17 557
rect 241 -619 275 557
rect 499 -619 533 557
rect 757 -619 791 557
rect 1015 -619 1049 557
rect 1273 -619 1307 557
rect 1531 -619 1565 557
<< mvpsubdiff >>
rect -1711 779 1711 791
rect -1711 745 -1603 779
rect 1603 745 1711 779
rect -1711 733 1711 745
rect -1711 546 -1653 733
rect -1711 -546 -1699 546
rect -1665 -546 -1653 546
rect -1711 -733 -1653 -546
rect 1653 546 1711 733
rect 1653 -546 1665 546
rect 1699 -546 1711 546
rect 1653 -733 1711 -546
rect -1711 -745 1711 -733
rect -1711 -779 -1603 -745
rect 1603 -779 1711 -745
rect -1711 -791 1711 -779
<< mvpsubdiffcont >>
rect -1603 745 1603 779
rect -1699 -546 -1665 546
rect 1665 -546 1699 546
rect -1603 -779 1603 -745
<< poly >>
rect -1502 641 -1336 657
rect -1502 624 -1486 641
rect -1519 607 -1486 624
rect -1352 624 -1336 641
rect -1244 641 -1078 657
rect -1244 624 -1228 641
rect -1352 607 -1319 624
rect -1519 569 -1319 607
rect -1261 607 -1228 624
rect -1094 624 -1078 641
rect -986 641 -820 657
rect -986 624 -970 641
rect -1094 607 -1061 624
rect -1261 569 -1061 607
rect -1003 607 -970 624
rect -836 624 -820 641
rect -728 641 -562 657
rect -728 624 -712 641
rect -836 607 -803 624
rect -1003 569 -803 607
rect -745 607 -712 624
rect -578 624 -562 641
rect -470 641 -304 657
rect -470 624 -454 641
rect -578 607 -545 624
rect -745 569 -545 607
rect -487 607 -454 624
rect -320 624 -304 641
rect -212 641 -46 657
rect -212 624 -196 641
rect -320 607 -287 624
rect -487 569 -287 607
rect -229 607 -196 624
rect -62 624 -46 641
rect 46 641 212 657
rect 46 624 62 641
rect -62 607 -29 624
rect -229 569 -29 607
rect 29 607 62 624
rect 196 624 212 641
rect 304 641 470 657
rect 304 624 320 641
rect 196 607 229 624
rect 29 569 229 607
rect 287 607 320 624
rect 454 624 470 641
rect 562 641 728 657
rect 562 624 578 641
rect 454 607 487 624
rect 287 569 487 607
rect 545 607 578 624
rect 712 624 728 641
rect 820 641 986 657
rect 820 624 836 641
rect 712 607 745 624
rect 545 569 745 607
rect 803 607 836 624
rect 970 624 986 641
rect 1078 641 1244 657
rect 1078 624 1094 641
rect 970 607 1003 624
rect 803 569 1003 607
rect 1061 607 1094 624
rect 1228 624 1244 641
rect 1336 641 1502 657
rect 1336 624 1352 641
rect 1228 607 1261 624
rect 1061 569 1261 607
rect 1319 607 1352 624
rect 1486 624 1502 641
rect 1486 607 1519 624
rect 1319 569 1519 607
rect -1519 -657 -1319 -631
rect -1261 -657 -1061 -631
rect -1003 -657 -803 -631
rect -745 -657 -545 -631
rect -487 -657 -287 -631
rect -229 -657 -29 -631
rect 29 -657 229 -631
rect 287 -657 487 -631
rect 545 -657 745 -631
rect 803 -657 1003 -631
rect 1061 -657 1261 -631
rect 1319 -657 1519 -631
<< polycont >>
rect -1486 607 -1352 641
rect -1228 607 -1094 641
rect -970 607 -836 641
rect -712 607 -578 641
rect -454 607 -320 641
rect -196 607 -62 641
rect 62 607 196 641
rect 320 607 454 641
rect 578 607 712 641
rect 836 607 970 641
rect 1094 607 1228 641
rect 1352 607 1486 641
<< locali >>
rect -1699 745 -1603 779
rect 1603 745 1699 779
rect -1699 546 -1665 745
rect -1699 -745 -1665 -546
rect -1565 557 -1531 573
rect -1565 -635 -1531 -619
rect -1307 557 -1273 573
rect -1307 -635 -1273 -619
rect -1049 557 -1015 573
rect -1049 -635 -1015 -619
rect -791 557 -757 573
rect -791 -635 -757 -619
rect -533 557 -499 573
rect -533 -635 -499 -619
rect -275 557 -241 573
rect -275 -635 -241 -619
rect -17 557 17 573
rect -17 -635 17 -619
rect 241 557 275 573
rect 241 -635 275 -619
rect 499 557 533 573
rect 499 -635 533 -619
rect 757 557 791 573
rect 757 -635 791 -619
rect 1015 557 1049 573
rect 1015 -635 1049 -619
rect 1273 557 1307 573
rect 1273 -635 1307 -619
rect 1531 557 1565 573
rect 1531 -635 1565 -619
rect 1665 546 1699 745
rect 1665 -745 1699 -546
rect -1699 -779 -1603 -745
rect 1603 -779 1699 -745
<< viali >>
rect -1503 607 -1486 641
rect -1486 607 -1352 641
rect -1352 607 -1335 641
rect -1245 607 -1228 641
rect -1228 607 -1094 641
rect -1094 607 -1077 641
rect -987 607 -970 641
rect -970 607 -836 641
rect -836 607 -819 641
rect -729 607 -712 641
rect -712 607 -578 641
rect -578 607 -561 641
rect -471 607 -454 641
rect -454 607 -320 641
rect -320 607 -303 641
rect -213 607 -196 641
rect -196 607 -62 641
rect -62 607 -45 641
rect 45 607 62 641
rect 62 607 196 641
rect 196 607 213 641
rect 303 607 320 641
rect 320 607 454 641
rect 454 607 471 641
rect 561 607 578 641
rect 578 607 712 641
rect 712 607 729 641
rect 819 607 836 641
rect 836 607 970 641
rect 970 607 987 641
rect 1077 607 1094 641
rect 1094 607 1228 641
rect 1228 607 1245 641
rect 1335 607 1352 641
rect 1352 607 1486 641
rect 1486 607 1503 641
rect -1565 -619 -1531 557
rect -1307 -619 -1273 557
rect -1049 -619 -1015 557
rect -791 -619 -757 557
rect -533 -619 -499 557
rect -275 -619 -241 557
rect -17 -619 17 557
rect 241 -619 275 557
rect 499 -619 533 557
rect 757 -619 791 557
rect 1015 -619 1049 557
rect 1273 -619 1307 557
rect 1531 -619 1565 557
<< metal1 >>
rect -1515 641 -1323 647
rect -1515 607 -1503 641
rect -1335 607 -1323 641
rect -1515 601 -1323 607
rect -1257 641 -1065 647
rect -1257 607 -1245 641
rect -1077 607 -1065 641
rect -1257 601 -1065 607
rect -999 641 -807 647
rect -999 607 -987 641
rect -819 607 -807 641
rect -999 601 -807 607
rect -741 641 -549 647
rect -741 607 -729 641
rect -561 607 -549 641
rect -741 601 -549 607
rect -483 641 -291 647
rect -483 607 -471 641
rect -303 607 -291 641
rect -483 601 -291 607
rect -225 641 -33 647
rect -225 607 -213 641
rect -45 607 -33 641
rect -225 601 -33 607
rect 33 641 225 647
rect 33 607 45 641
rect 213 607 225 641
rect 33 601 225 607
rect 291 641 483 647
rect 291 607 303 641
rect 471 607 483 641
rect 291 601 483 607
rect 549 641 741 647
rect 549 607 561 641
rect 729 607 741 641
rect 549 601 741 607
rect 807 641 999 647
rect 807 607 819 641
rect 987 607 999 641
rect 807 601 999 607
rect 1065 641 1257 647
rect 1065 607 1077 641
rect 1245 607 1257 641
rect 1065 601 1257 607
rect 1323 641 1515 647
rect 1323 607 1335 641
rect 1503 607 1515 641
rect 1323 601 1515 607
rect -1571 557 -1525 569
rect -1571 -619 -1565 557
rect -1531 -619 -1525 557
rect -1571 -631 -1525 -619
rect -1313 557 -1267 569
rect -1313 -619 -1307 557
rect -1273 -619 -1267 557
rect -1313 -631 -1267 -619
rect -1055 557 -1009 569
rect -1055 -619 -1049 557
rect -1015 -619 -1009 557
rect -1055 -631 -1009 -619
rect -797 557 -751 569
rect -797 -619 -791 557
rect -757 -619 -751 557
rect -797 -631 -751 -619
rect -539 557 -493 569
rect -539 -619 -533 557
rect -499 -619 -493 557
rect -539 -631 -493 -619
rect -281 557 -235 569
rect -281 -619 -275 557
rect -241 -619 -235 557
rect -281 -631 -235 -619
rect -23 557 23 569
rect -23 -619 -17 557
rect 17 -619 23 557
rect -23 -631 23 -619
rect 235 557 281 569
rect 235 -619 241 557
rect 275 -619 281 557
rect 235 -631 281 -619
rect 493 557 539 569
rect 493 -619 499 557
rect 533 -619 539 557
rect 493 -631 539 -619
rect 751 557 797 569
rect 751 -619 757 557
rect 791 -619 797 557
rect 751 -631 797 -619
rect 1009 557 1055 569
rect 1009 -619 1015 557
rect 1049 -619 1055 557
rect 1009 -631 1055 -619
rect 1267 557 1313 569
rect 1267 -619 1273 557
rect 1307 -619 1313 557
rect 1267 -631 1313 -619
rect 1525 557 1571 569
rect 1525 -619 1531 557
rect 1565 -619 1571 557
rect 1525 -631 1571 -619
<< properties >>
string FIXED_BBOX -1682 -762 1682 762
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 6 l 1 m 1 nf 12 diffcov 100 polycov 80 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 80 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
