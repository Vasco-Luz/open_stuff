magic
tech sky130A
timestamp 1693418132
<< pwell >>
rect -443 -229 443 229
<< mvnmos >>
rect -329 -100 -129 100
rect -100 -100 100 100
rect 129 -100 329 100
<< mvndiff >>
rect -358 94 -329 100
rect -358 -94 -352 94
rect -335 -94 -329 94
rect -358 -100 -329 -94
rect -129 94 -100 100
rect -129 -94 -123 94
rect -106 -94 -100 94
rect -129 -100 -100 -94
rect 100 94 129 100
rect 100 -94 106 94
rect 123 -94 129 94
rect 100 -100 129 -94
rect 329 94 358 100
rect 329 -94 335 94
rect 352 -94 358 94
rect 329 -100 358 -94
<< mvndiffc >>
rect -352 -94 -335 94
rect -123 -94 -106 94
rect 106 -94 123 94
rect 335 -94 352 94
<< mvpsubdiff >>
rect -425 205 425 211
rect -425 188 -371 205
rect 371 188 425 205
rect -425 182 425 188
rect -425 157 -396 182
rect -425 -157 -419 157
rect -402 -157 -396 157
rect 396 157 425 182
rect -425 -182 -396 -157
rect 396 -157 402 157
rect 419 -157 425 157
rect 396 -182 425 -157
rect -425 -188 425 -182
rect -425 -205 -371 -188
rect 371 -205 425 -188
rect -425 -211 425 -205
<< mvpsubdiffcont >>
rect -371 188 371 205
rect -419 -157 -402 157
rect 402 -157 419 157
rect -371 -205 371 -188
<< poly >>
rect -329 136 -129 144
rect -329 119 -321 136
rect -137 119 -129 136
rect -329 100 -129 119
rect -100 136 100 144
rect -100 119 -92 136
rect 92 119 100 136
rect -100 100 100 119
rect 129 136 329 144
rect 129 119 137 136
rect 321 119 329 136
rect 129 100 329 119
rect -329 -119 -129 -100
rect -329 -136 -321 -119
rect -137 -136 -129 -119
rect -329 -144 -129 -136
rect -100 -119 100 -100
rect -100 -136 -92 -119
rect 92 -136 100 -119
rect -100 -144 100 -136
rect 129 -119 329 -100
rect 129 -136 137 -119
rect 321 -136 329 -119
rect 129 -144 329 -136
<< polycont >>
rect -321 119 -137 136
rect -92 119 92 136
rect 137 119 321 136
rect -321 -136 -137 -119
rect -92 -136 92 -119
rect 137 -136 321 -119
<< locali >>
rect -419 188 -371 205
rect 371 188 419 205
rect -419 157 -402 188
rect 402 157 419 188
rect -329 119 -321 136
rect -137 119 -129 136
rect -100 119 -92 136
rect 92 119 100 136
rect 129 119 137 136
rect 321 119 329 136
rect -352 94 -335 102
rect -352 -102 -335 -94
rect -123 94 -106 102
rect -123 -102 -106 -94
rect 106 94 123 102
rect 106 -102 123 -94
rect 335 94 352 102
rect 335 -102 352 -94
rect -329 -136 -321 -119
rect -137 -136 -129 -119
rect -100 -136 -92 -119
rect 92 -136 100 -119
rect 129 -136 137 -119
rect 321 -136 329 -119
rect -419 -188 -402 -157
rect 402 -188 419 -157
rect -419 -205 -371 -188
rect 371 -205 419 -188
<< viali >>
rect -321 119 -137 136
rect -92 119 92 136
rect 137 119 321 136
rect -352 -94 -335 94
rect -123 -94 -106 94
rect 106 -94 123 94
rect 335 -94 352 94
rect -321 -136 -137 -119
rect -92 -136 92 -119
rect 137 -136 321 -119
<< metal1 >>
rect -327 136 -131 139
rect -327 119 -321 136
rect -137 119 -131 136
rect -327 116 -131 119
rect -98 136 98 139
rect -98 119 -92 136
rect 92 119 98 136
rect -98 116 98 119
rect 131 136 327 139
rect 131 119 137 136
rect 321 119 327 136
rect 131 116 327 119
rect -355 94 -332 100
rect -355 -94 -352 94
rect -335 -94 -332 94
rect -355 -100 -332 -94
rect -126 94 -103 100
rect -126 -94 -123 94
rect -106 -94 -103 94
rect -126 -100 -103 -94
rect 103 94 126 100
rect 103 -94 106 94
rect 123 -94 126 94
rect 103 -100 126 -94
rect 332 94 355 100
rect 332 -94 335 94
rect 352 -94 355 94
rect 332 -100 355 -94
rect -327 -119 -131 -116
rect -327 -136 -321 -119
rect -137 -136 -131 -119
rect -327 -139 -131 -136
rect -98 -119 98 -116
rect -98 -136 -92 -119
rect 92 -136 98 -119
rect -98 -139 98 -136
rect 131 -119 327 -116
rect 131 -136 137 -119
rect 321 -136 327 -119
rect 131 -139 327 -136
<< properties >>
string FIXED_BBOX -410 -196 410 196
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 2 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
