magic
tech sky130A
magscale 1 2
timestamp 1693011900
<< pwell >>
rect -352 -798 352 798
<< psubdiff >>
rect -316 728 -220 762
rect 220 728 316 762
rect -316 666 -282 728
rect 282 666 316 728
rect -316 -728 -282 -666
rect 282 -728 316 -666
rect -316 -762 -220 -728
rect 220 -762 316 -728
<< psubdiffcont >>
rect -220 728 220 762
rect -316 -666 -282 666
rect 282 -666 316 666
rect -220 -762 220 -728
<< xpolycontact >>
rect -186 200 -48 632
rect -186 -632 -48 -200
rect 48 200 186 632
rect 48 -632 186 -200
<< ppolyres >>
rect -186 -200 -48 200
rect 48 -200 186 200
<< locali >>
rect -316 728 -220 762
rect 220 728 316 762
rect -316 666 -282 728
rect 282 666 316 728
rect -316 -728 -282 -666
rect 282 -728 316 -666
rect -316 -762 -220 -728
rect 220 -762 316 -728
<< viali >>
rect -170 217 -64 614
rect 64 217 170 614
rect -170 -614 -64 -217
rect 64 -614 170 -217
<< metal1 >>
rect -176 614 -58 626
rect -176 217 -170 614
rect -64 217 -58 614
rect -176 205 -58 217
rect 58 614 176 626
rect 58 217 64 614
rect 170 217 176 614
rect 58 205 176 217
rect -176 -217 -58 -205
rect -176 -614 -170 -217
rect -64 -614 -58 -217
rect -176 -626 -58 -614
rect 58 -217 176 -205
rect 58 -614 64 -217
rect 170 -614 176 -217
rect 58 -626 176 -614
<< properties >>
string FIXED_BBOX -299 -745 299 745
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.69 l 2 m 1 nx 2 wmin 0.690 lmin 0.50 rho 319.8 val 1.491k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
