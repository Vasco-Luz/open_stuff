magic
tech sky130A
magscale 1 2
timestamp 1693418132
<< pwell >>
rect -1344 -427 1344 427
<< mvnmos >>
rect -1116 -231 -716 169
rect -658 -231 -258 169
rect -200 -231 200 169
rect 258 -231 658 169
rect 716 -231 1116 169
<< mvndiff >>
rect -1174 157 -1116 169
rect -1174 -219 -1162 157
rect -1128 -219 -1116 157
rect -1174 -231 -1116 -219
rect -716 157 -658 169
rect -716 -219 -704 157
rect -670 -219 -658 157
rect -716 -231 -658 -219
rect -258 157 -200 169
rect -258 -219 -246 157
rect -212 -219 -200 157
rect -258 -231 -200 -219
rect 200 157 258 169
rect 200 -219 212 157
rect 246 -219 258 157
rect 200 -231 258 -219
rect 658 157 716 169
rect 658 -219 670 157
rect 704 -219 716 157
rect 658 -231 716 -219
rect 1116 157 1174 169
rect 1116 -219 1128 157
rect 1162 -219 1174 157
rect 1116 -231 1174 -219
<< mvndiffc >>
rect -1162 -219 -1128 157
rect -704 -219 -670 157
rect -246 -219 -212 157
rect 212 -219 246 157
rect 670 -219 704 157
rect 1128 -219 1162 157
<< mvpsubdiff >>
rect -1308 379 1308 391
rect -1308 345 -1200 379
rect 1200 345 1308 379
rect -1308 333 1308 345
rect -1308 283 -1250 333
rect -1308 -283 -1296 283
rect -1262 -283 -1250 283
rect 1250 283 1308 333
rect -1308 -333 -1250 -283
rect 1250 -283 1262 283
rect 1296 -283 1308 283
rect 1250 -333 1308 -283
rect -1308 -345 1308 -333
rect -1308 -379 -1200 -345
rect 1200 -379 1308 -345
rect -1308 -391 1308 -379
<< mvpsubdiffcont >>
rect -1200 345 1200 379
rect -1296 -283 -1262 283
rect 1262 -283 1296 283
rect -1200 -379 1200 -345
<< poly >>
rect -1024 241 -808 257
rect -1024 224 -1008 241
rect -1116 207 -1008 224
rect -824 224 -808 241
rect -566 241 -350 257
rect -566 224 -550 241
rect -824 207 -716 224
rect -1116 169 -716 207
rect -658 207 -550 224
rect -366 224 -350 241
rect -108 241 108 257
rect -108 224 -92 241
rect -366 207 -258 224
rect -658 169 -258 207
rect -200 207 -92 224
rect 92 224 108 241
rect 350 241 566 257
rect 350 224 366 241
rect 92 207 200 224
rect -200 169 200 207
rect 258 207 366 224
rect 550 224 566 241
rect 808 241 1024 257
rect 808 224 824 241
rect 550 207 658 224
rect 258 169 658 207
rect 716 207 824 224
rect 1008 224 1024 241
rect 1008 207 1116 224
rect 716 169 1116 207
rect -1116 -257 -716 -231
rect -658 -257 -258 -231
rect -200 -257 200 -231
rect 258 -257 658 -231
rect 716 -257 1116 -231
<< polycont >>
rect -1008 207 -824 241
rect -550 207 -366 241
rect -92 207 92 241
rect 366 207 550 241
rect 824 207 1008 241
<< locali >>
rect -1296 345 -1200 379
rect 1200 345 1296 379
rect -1296 283 -1262 345
rect 1262 283 1296 345
rect -1024 207 -1008 241
rect -824 207 -808 241
rect -566 207 -550 241
rect -366 207 -350 241
rect -108 207 -92 241
rect 92 207 108 241
rect 350 207 366 241
rect 550 207 566 241
rect 808 207 824 241
rect 1008 207 1024 241
rect -1162 157 -1128 173
rect -1162 -235 -1128 -219
rect -704 157 -670 173
rect -704 -235 -670 -219
rect -246 157 -212 173
rect -246 -235 -212 -219
rect 212 157 246 173
rect 212 -235 246 -219
rect 670 157 704 173
rect 670 -235 704 -219
rect 1128 157 1162 173
rect 1128 -235 1162 -219
rect -1296 -345 -1262 -283
rect 1262 -345 1296 -283
rect -1296 -379 -1200 -345
rect 1200 -379 1296 -345
<< viali >>
rect -1008 207 -824 241
rect -550 207 -366 241
rect -92 207 92 241
rect 366 207 550 241
rect 824 207 1008 241
rect -1162 -200 -1128 138
rect -704 -200 -670 138
rect -246 -200 -212 138
rect 212 -200 246 138
rect 670 -200 704 138
rect 1128 -200 1162 138
<< metal1 >>
rect -1020 241 -812 247
rect -1020 207 -1008 241
rect -824 207 -812 241
rect -1020 201 -812 207
rect -562 241 -354 247
rect -562 207 -550 241
rect -366 207 -354 241
rect -562 201 -354 207
rect -104 241 104 247
rect -104 207 -92 241
rect 92 207 104 241
rect -104 201 104 207
rect 354 241 562 247
rect 354 207 366 241
rect 550 207 562 241
rect 354 201 562 207
rect 812 241 1020 247
rect 812 207 824 241
rect 1008 207 1020 241
rect 812 201 1020 207
rect -1168 138 -1122 150
rect -1168 -200 -1162 138
rect -1128 -200 -1122 138
rect -1168 -212 -1122 -200
rect -710 138 -664 150
rect -710 -200 -704 138
rect -670 -200 -664 138
rect -710 -212 -664 -200
rect -252 138 -206 150
rect -252 -200 -246 138
rect -212 -200 -206 138
rect -252 -212 -206 -200
rect 206 138 252 150
rect 206 -200 212 138
rect 246 -200 252 138
rect 206 -212 252 -200
rect 664 138 710 150
rect 664 -200 670 138
rect 704 -200 710 138
rect 664 -212 710 -200
rect 1122 138 1168 150
rect 1122 -200 1128 138
rect 1162 -200 1168 138
rect 1122 -212 1168 -200
<< properties >>
string FIXED_BBOX -1279 -362 1279 362
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 2 m 1 nf 5 diffcov 100 polycov 50 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 90 viadrn 90 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
