magic
tech sky130A
magscale 1 2
timestamp 1693420066
<< error_p >>
rect -1530 541 -1472 547
rect -1372 541 -1314 547
rect -1214 541 -1156 547
rect -1056 541 -998 547
rect -898 541 -840 547
rect -740 541 -682 547
rect -582 541 -524 547
rect -424 541 -366 547
rect -266 541 -208 547
rect -108 541 -50 547
rect 50 541 108 547
rect 208 541 266 547
rect 366 541 424 547
rect 524 541 582 547
rect 682 541 740 547
rect 840 541 898 547
rect 998 541 1056 547
rect 1156 541 1214 547
rect 1314 541 1372 547
rect 1472 541 1530 547
rect -1530 507 -1518 541
rect -1372 507 -1360 541
rect -1214 507 -1202 541
rect -1056 507 -1044 541
rect -898 507 -886 541
rect -740 507 -728 541
rect -582 507 -570 541
rect -424 507 -412 541
rect -266 507 -254 541
rect -108 507 -96 541
rect 50 507 62 541
rect 208 507 220 541
rect 366 507 378 541
rect 524 507 536 541
rect 682 507 694 541
rect 840 507 852 541
rect 998 507 1010 541
rect 1156 507 1168 541
rect 1314 507 1326 541
rect 1472 507 1484 541
rect -1530 501 -1472 507
rect -1372 501 -1314 507
rect -1214 501 -1156 507
rect -1056 501 -998 507
rect -898 501 -840 507
rect -740 501 -682 507
rect -582 501 -524 507
rect -424 501 -366 507
rect -266 501 -208 507
rect -108 501 -50 507
rect 50 501 108 507
rect 208 501 266 507
rect 366 501 424 507
rect 524 501 582 507
rect 682 501 740 507
rect 840 501 898 507
rect 998 501 1056 507
rect 1156 501 1214 507
rect 1314 501 1372 507
rect 1472 501 1530 507
<< pwell >>
rect -1779 -727 1779 727
<< mvnmos >>
rect -1551 -531 -1451 469
rect -1393 -531 -1293 469
rect -1235 -531 -1135 469
rect -1077 -531 -977 469
rect -919 -531 -819 469
rect -761 -531 -661 469
rect -603 -531 -503 469
rect -445 -531 -345 469
rect -287 -531 -187 469
rect -129 -531 -29 469
rect 29 -531 129 469
rect 187 -531 287 469
rect 345 -531 445 469
rect 503 -531 603 469
rect 661 -531 761 469
rect 819 -531 919 469
rect 977 -531 1077 469
rect 1135 -531 1235 469
rect 1293 -531 1393 469
rect 1451 -531 1551 469
<< mvndiff >>
rect -1609 457 -1551 469
rect -1609 -519 -1597 457
rect -1563 -519 -1551 457
rect -1609 -531 -1551 -519
rect -1451 457 -1393 469
rect -1451 -519 -1439 457
rect -1405 -519 -1393 457
rect -1451 -531 -1393 -519
rect -1293 457 -1235 469
rect -1293 -519 -1281 457
rect -1247 -519 -1235 457
rect -1293 -531 -1235 -519
rect -1135 457 -1077 469
rect -1135 -519 -1123 457
rect -1089 -519 -1077 457
rect -1135 -531 -1077 -519
rect -977 457 -919 469
rect -977 -519 -965 457
rect -931 -519 -919 457
rect -977 -531 -919 -519
rect -819 457 -761 469
rect -819 -519 -807 457
rect -773 -519 -761 457
rect -819 -531 -761 -519
rect -661 457 -603 469
rect -661 -519 -649 457
rect -615 -519 -603 457
rect -661 -531 -603 -519
rect -503 457 -445 469
rect -503 -519 -491 457
rect -457 -519 -445 457
rect -503 -531 -445 -519
rect -345 457 -287 469
rect -345 -519 -333 457
rect -299 -519 -287 457
rect -345 -531 -287 -519
rect -187 457 -129 469
rect -187 -519 -175 457
rect -141 -519 -129 457
rect -187 -531 -129 -519
rect -29 457 29 469
rect -29 -519 -17 457
rect 17 -519 29 457
rect -29 -531 29 -519
rect 129 457 187 469
rect 129 -519 141 457
rect 175 -519 187 457
rect 129 -531 187 -519
rect 287 457 345 469
rect 287 -519 299 457
rect 333 -519 345 457
rect 287 -531 345 -519
rect 445 457 503 469
rect 445 -519 457 457
rect 491 -519 503 457
rect 445 -531 503 -519
rect 603 457 661 469
rect 603 -519 615 457
rect 649 -519 661 457
rect 603 -531 661 -519
rect 761 457 819 469
rect 761 -519 773 457
rect 807 -519 819 457
rect 761 -531 819 -519
rect 919 457 977 469
rect 919 -519 931 457
rect 965 -519 977 457
rect 919 -531 977 -519
rect 1077 457 1135 469
rect 1077 -519 1089 457
rect 1123 -519 1135 457
rect 1077 -531 1135 -519
rect 1235 457 1293 469
rect 1235 -519 1247 457
rect 1281 -519 1293 457
rect 1235 -531 1293 -519
rect 1393 457 1451 469
rect 1393 -519 1405 457
rect 1439 -519 1451 457
rect 1393 -531 1451 -519
rect 1551 457 1609 469
rect 1551 -519 1563 457
rect 1597 -519 1609 457
rect 1551 -531 1609 -519
<< mvndiffc >>
rect -1597 -519 -1563 457
rect -1439 -519 -1405 457
rect -1281 -519 -1247 457
rect -1123 -519 -1089 457
rect -965 -519 -931 457
rect -807 -519 -773 457
rect -649 -519 -615 457
rect -491 -519 -457 457
rect -333 -519 -299 457
rect -175 -519 -141 457
rect -17 -519 17 457
rect 141 -519 175 457
rect 299 -519 333 457
rect 457 -519 491 457
rect 615 -519 649 457
rect 773 -519 807 457
rect 931 -519 965 457
rect 1089 -519 1123 457
rect 1247 -519 1281 457
rect 1405 -519 1439 457
rect 1563 -519 1597 457
<< mvpsubdiff >>
rect -1743 679 1743 691
rect -1743 645 -1635 679
rect 1635 645 1743 679
rect -1743 633 1743 645
rect -1743 583 -1685 633
rect -1743 -583 -1731 583
rect -1697 -583 -1685 583
rect 1685 583 1743 633
rect -1743 -633 -1685 -583
rect 1685 -583 1697 583
rect 1731 -583 1743 583
rect 1685 -633 1743 -583
rect -1743 -645 1743 -633
rect -1743 -679 -1635 -645
rect 1635 -679 1743 -645
rect -1743 -691 1743 -679
<< mvpsubdiffcont >>
rect -1635 645 1635 679
rect -1731 -583 -1697 583
rect 1697 -583 1731 583
rect -1635 -679 1635 -645
<< poly >>
rect -1534 541 -1468 557
rect -1534 524 -1518 541
rect -1551 507 -1518 524
rect -1484 524 -1468 541
rect -1376 541 -1310 557
rect -1376 524 -1360 541
rect -1484 507 -1451 524
rect -1551 469 -1451 507
rect -1393 507 -1360 524
rect -1326 524 -1310 541
rect -1218 541 -1152 557
rect -1218 524 -1202 541
rect -1326 507 -1293 524
rect -1393 469 -1293 507
rect -1235 507 -1202 524
rect -1168 524 -1152 541
rect -1060 541 -994 557
rect -1060 524 -1044 541
rect -1168 507 -1135 524
rect -1235 469 -1135 507
rect -1077 507 -1044 524
rect -1010 524 -994 541
rect -902 541 -836 557
rect -902 524 -886 541
rect -1010 507 -977 524
rect -1077 469 -977 507
rect -919 507 -886 524
rect -852 524 -836 541
rect -744 541 -678 557
rect -744 524 -728 541
rect -852 507 -819 524
rect -919 469 -819 507
rect -761 507 -728 524
rect -694 524 -678 541
rect -586 541 -520 557
rect -586 524 -570 541
rect -694 507 -661 524
rect -761 469 -661 507
rect -603 507 -570 524
rect -536 524 -520 541
rect -428 541 -362 557
rect -428 524 -412 541
rect -536 507 -503 524
rect -603 469 -503 507
rect -445 507 -412 524
rect -378 524 -362 541
rect -270 541 -204 557
rect -270 524 -254 541
rect -378 507 -345 524
rect -445 469 -345 507
rect -287 507 -254 524
rect -220 524 -204 541
rect -112 541 -46 557
rect -112 524 -96 541
rect -220 507 -187 524
rect -287 469 -187 507
rect -129 507 -96 524
rect -62 524 -46 541
rect 46 541 112 557
rect 46 524 62 541
rect -62 507 -29 524
rect -129 469 -29 507
rect 29 507 62 524
rect 96 524 112 541
rect 204 541 270 557
rect 204 524 220 541
rect 96 507 129 524
rect 29 469 129 507
rect 187 507 220 524
rect 254 524 270 541
rect 362 541 428 557
rect 362 524 378 541
rect 254 507 287 524
rect 187 469 287 507
rect 345 507 378 524
rect 412 524 428 541
rect 520 541 586 557
rect 520 524 536 541
rect 412 507 445 524
rect 345 469 445 507
rect 503 507 536 524
rect 570 524 586 541
rect 678 541 744 557
rect 678 524 694 541
rect 570 507 603 524
rect 503 469 603 507
rect 661 507 694 524
rect 728 524 744 541
rect 836 541 902 557
rect 836 524 852 541
rect 728 507 761 524
rect 661 469 761 507
rect 819 507 852 524
rect 886 524 902 541
rect 994 541 1060 557
rect 994 524 1010 541
rect 886 507 919 524
rect 819 469 919 507
rect 977 507 1010 524
rect 1044 524 1060 541
rect 1152 541 1218 557
rect 1152 524 1168 541
rect 1044 507 1077 524
rect 977 469 1077 507
rect 1135 507 1168 524
rect 1202 524 1218 541
rect 1310 541 1376 557
rect 1310 524 1326 541
rect 1202 507 1235 524
rect 1135 469 1235 507
rect 1293 507 1326 524
rect 1360 524 1376 541
rect 1468 541 1534 557
rect 1468 524 1484 541
rect 1360 507 1393 524
rect 1293 469 1393 507
rect 1451 507 1484 524
rect 1518 524 1534 541
rect 1518 507 1551 524
rect 1451 469 1551 507
rect -1551 -557 -1451 -531
rect -1393 -557 -1293 -531
rect -1235 -557 -1135 -531
rect -1077 -557 -977 -531
rect -919 -557 -819 -531
rect -761 -557 -661 -531
rect -603 -557 -503 -531
rect -445 -557 -345 -531
rect -287 -557 -187 -531
rect -129 -557 -29 -531
rect 29 -557 129 -531
rect 187 -557 287 -531
rect 345 -557 445 -531
rect 503 -557 603 -531
rect 661 -557 761 -531
rect 819 -557 919 -531
rect 977 -557 1077 -531
rect 1135 -557 1235 -531
rect 1293 -557 1393 -531
rect 1451 -557 1551 -531
<< polycont >>
rect -1518 507 -1484 541
rect -1360 507 -1326 541
rect -1202 507 -1168 541
rect -1044 507 -1010 541
rect -886 507 -852 541
rect -728 507 -694 541
rect -570 507 -536 541
rect -412 507 -378 541
rect -254 507 -220 541
rect -96 507 -62 541
rect 62 507 96 541
rect 220 507 254 541
rect 378 507 412 541
rect 536 507 570 541
rect 694 507 728 541
rect 852 507 886 541
rect 1010 507 1044 541
rect 1168 507 1202 541
rect 1326 507 1360 541
rect 1484 507 1518 541
<< locali >>
rect -1731 645 -1635 679
rect 1635 645 1731 679
rect -1731 583 -1697 645
rect 1697 583 1731 645
rect -1534 507 -1518 541
rect -1484 507 -1468 541
rect -1376 507 -1360 541
rect -1326 507 -1310 541
rect -1218 507 -1202 541
rect -1168 507 -1152 541
rect -1060 507 -1044 541
rect -1010 507 -994 541
rect -902 507 -886 541
rect -852 507 -836 541
rect -744 507 -728 541
rect -694 507 -678 541
rect -586 507 -570 541
rect -536 507 -520 541
rect -428 507 -412 541
rect -378 507 -362 541
rect -270 507 -254 541
rect -220 507 -204 541
rect -112 507 -96 541
rect -62 507 -46 541
rect 46 507 62 541
rect 96 507 112 541
rect 204 507 220 541
rect 254 507 270 541
rect 362 507 378 541
rect 412 507 428 541
rect 520 507 536 541
rect 570 507 586 541
rect 678 507 694 541
rect 728 507 744 541
rect 836 507 852 541
rect 886 507 902 541
rect 994 507 1010 541
rect 1044 507 1060 541
rect 1152 507 1168 541
rect 1202 507 1218 541
rect 1310 507 1326 541
rect 1360 507 1376 541
rect 1468 507 1484 541
rect 1518 507 1534 541
rect -1597 457 -1563 473
rect -1597 -535 -1563 -519
rect -1439 457 -1405 473
rect -1439 -535 -1405 -519
rect -1281 457 -1247 473
rect -1281 -535 -1247 -519
rect -1123 457 -1089 473
rect -1123 -535 -1089 -519
rect -965 457 -931 473
rect -965 -535 -931 -519
rect -807 457 -773 473
rect -807 -535 -773 -519
rect -649 457 -615 473
rect -649 -535 -615 -519
rect -491 457 -457 473
rect -491 -535 -457 -519
rect -333 457 -299 473
rect -333 -535 -299 -519
rect -175 457 -141 473
rect -175 -535 -141 -519
rect -17 457 17 473
rect -17 -535 17 -519
rect 141 457 175 473
rect 141 -535 175 -519
rect 299 457 333 473
rect 299 -535 333 -519
rect 457 457 491 473
rect 457 -535 491 -519
rect 615 457 649 473
rect 615 -535 649 -519
rect 773 457 807 473
rect 773 -535 807 -519
rect 931 457 965 473
rect 931 -535 965 -519
rect 1089 457 1123 473
rect 1089 -535 1123 -519
rect 1247 457 1281 473
rect 1247 -535 1281 -519
rect 1405 457 1439 473
rect 1405 -535 1439 -519
rect 1563 457 1597 473
rect 1563 -535 1597 -519
rect -1731 -645 -1697 -583
rect 1697 -645 1731 -583
rect -1731 -679 -1635 -645
rect 1635 -679 1731 -645
<< viali >>
rect -1518 507 -1484 541
rect -1360 507 -1326 541
rect -1202 507 -1168 541
rect -1044 507 -1010 541
rect -886 507 -852 541
rect -728 507 -694 541
rect -570 507 -536 541
rect -412 507 -378 541
rect -254 507 -220 541
rect -96 507 -62 541
rect 62 507 96 541
rect 220 507 254 541
rect 378 507 412 541
rect 536 507 570 541
rect 694 507 728 541
rect 852 507 886 541
rect 1010 507 1044 541
rect 1168 507 1202 541
rect 1326 507 1360 541
rect 1484 507 1518 541
rect -1597 -519 -1563 457
rect -1439 -519 -1405 457
rect -1281 -519 -1247 457
rect -1123 -519 -1089 457
rect -965 -519 -931 457
rect -807 -519 -773 457
rect -649 -519 -615 457
rect -491 -519 -457 457
rect -333 -519 -299 457
rect -175 -519 -141 457
rect -17 -519 17 457
rect 141 -519 175 457
rect 299 -519 333 457
rect 457 -519 491 457
rect 615 -519 649 457
rect 773 -519 807 457
rect 931 -519 965 457
rect 1089 -519 1123 457
rect 1247 -519 1281 457
rect 1405 -519 1439 457
rect 1563 -519 1597 457
<< metal1 >>
rect -1530 541 -1472 547
rect -1530 507 -1518 541
rect -1484 507 -1472 541
rect -1530 501 -1472 507
rect -1372 541 -1314 547
rect -1372 507 -1360 541
rect -1326 507 -1314 541
rect -1372 501 -1314 507
rect -1214 541 -1156 547
rect -1214 507 -1202 541
rect -1168 507 -1156 541
rect -1214 501 -1156 507
rect -1056 541 -998 547
rect -1056 507 -1044 541
rect -1010 507 -998 541
rect -1056 501 -998 507
rect -898 541 -840 547
rect -898 507 -886 541
rect -852 507 -840 541
rect -898 501 -840 507
rect -740 541 -682 547
rect -740 507 -728 541
rect -694 507 -682 541
rect -740 501 -682 507
rect -582 541 -524 547
rect -582 507 -570 541
rect -536 507 -524 541
rect -582 501 -524 507
rect -424 541 -366 547
rect -424 507 -412 541
rect -378 507 -366 541
rect -424 501 -366 507
rect -266 541 -208 547
rect -266 507 -254 541
rect -220 507 -208 541
rect -266 501 -208 507
rect -108 541 -50 547
rect -108 507 -96 541
rect -62 507 -50 541
rect -108 501 -50 507
rect 50 541 108 547
rect 50 507 62 541
rect 96 507 108 541
rect 50 501 108 507
rect 208 541 266 547
rect 208 507 220 541
rect 254 507 266 541
rect 208 501 266 507
rect 366 541 424 547
rect 366 507 378 541
rect 412 507 424 541
rect 366 501 424 507
rect 524 541 582 547
rect 524 507 536 541
rect 570 507 582 541
rect 524 501 582 507
rect 682 541 740 547
rect 682 507 694 541
rect 728 507 740 541
rect 682 501 740 507
rect 840 541 898 547
rect 840 507 852 541
rect 886 507 898 541
rect 840 501 898 507
rect 998 541 1056 547
rect 998 507 1010 541
rect 1044 507 1056 541
rect 998 501 1056 507
rect 1156 541 1214 547
rect 1156 507 1168 541
rect 1202 507 1214 541
rect 1156 501 1214 507
rect 1314 541 1372 547
rect 1314 507 1326 541
rect 1360 507 1372 541
rect 1314 501 1372 507
rect 1472 541 1530 547
rect 1472 507 1484 541
rect 1518 507 1530 541
rect 1472 501 1530 507
rect -1603 457 -1557 469
rect -1603 -519 -1597 457
rect -1563 -519 -1557 457
rect -1603 -531 -1557 -519
rect -1445 457 -1399 469
rect -1445 -519 -1439 457
rect -1405 -519 -1399 457
rect -1445 -531 -1399 -519
rect -1287 457 -1241 469
rect -1287 -519 -1281 457
rect -1247 -519 -1241 457
rect -1287 -531 -1241 -519
rect -1129 457 -1083 469
rect -1129 -519 -1123 457
rect -1089 -519 -1083 457
rect -1129 -531 -1083 -519
rect -971 457 -925 469
rect -971 -519 -965 457
rect -931 -519 -925 457
rect -971 -531 -925 -519
rect -813 457 -767 469
rect -813 -519 -807 457
rect -773 -519 -767 457
rect -813 -531 -767 -519
rect -655 457 -609 469
rect -655 -519 -649 457
rect -615 -519 -609 457
rect -655 -531 -609 -519
rect -497 457 -451 469
rect -497 -519 -491 457
rect -457 -519 -451 457
rect -497 -531 -451 -519
rect -339 457 -293 469
rect -339 -519 -333 457
rect -299 -519 -293 457
rect -339 -531 -293 -519
rect -181 457 -135 469
rect -181 -519 -175 457
rect -141 -519 -135 457
rect -181 -531 -135 -519
rect -23 457 23 469
rect -23 -519 -17 457
rect 17 -519 23 457
rect -23 -531 23 -519
rect 135 457 181 469
rect 135 -519 141 457
rect 175 -519 181 457
rect 135 -531 181 -519
rect 293 457 339 469
rect 293 -519 299 457
rect 333 -519 339 457
rect 293 -531 339 -519
rect 451 457 497 469
rect 451 -519 457 457
rect 491 -519 497 457
rect 451 -531 497 -519
rect 609 457 655 469
rect 609 -519 615 457
rect 649 -519 655 457
rect 609 -531 655 -519
rect 767 457 813 469
rect 767 -519 773 457
rect 807 -519 813 457
rect 767 -531 813 -519
rect 925 457 971 469
rect 925 -519 931 457
rect 965 -519 971 457
rect 925 -531 971 -519
rect 1083 457 1129 469
rect 1083 -519 1089 457
rect 1123 -519 1129 457
rect 1083 -531 1129 -519
rect 1241 457 1287 469
rect 1241 -519 1247 457
rect 1281 -519 1287 457
rect 1241 -531 1287 -519
rect 1399 457 1445 469
rect 1399 -519 1405 457
rect 1439 -519 1445 457
rect 1399 -531 1445 -519
rect 1557 457 1603 469
rect 1557 -519 1563 457
rect 1597 -519 1603 457
rect 1557 -531 1603 -519
<< properties >>
string FIXED_BBOX -1714 -662 1714 662
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.5 m 1 nf 20 diffcov 100 polycov 50 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
