magic
tech sky130A
magscale 1 2
timestamp 1693050045
<< nwell >>
rect 332 122 420 130
<< poly >>
rect 561 -342 715 -326
rect 561 -376 571 -342
rect 705 -376 715 -342
rect 561 -388 715 -376
rect 819 -342 973 -326
rect 819 -376 829 -342
rect 963 -376 973 -342
rect 819 -388 973 -376
rect 1077 -342 1231 -326
rect 1077 -376 1087 -342
rect 1221 -376 1231 -342
rect 1077 -388 1231 -376
rect 1335 -342 1489 -326
rect 1335 -376 1345 -342
rect 1479 -376 1489 -342
rect 1335 -388 1489 -376
rect 1593 -342 1747 -326
rect 1593 -376 1603 -342
rect 1737 -376 1747 -342
rect 1593 -388 1747 -376
rect 1851 -342 2005 -326
rect 1851 -376 1861 -342
rect 1995 -376 2005 -342
rect 1851 -388 2005 -376
rect 2109 -342 2263 -326
rect 2109 -376 2119 -342
rect 2253 -376 2263 -342
rect 2109 -388 2263 -376
rect 2367 -342 2521 -326
rect 2367 -376 2377 -342
rect 2511 -376 2521 -342
rect 2367 -388 2521 -376
rect 2625 -342 2779 -326
rect 2625 -376 2635 -342
rect 2769 -376 2779 -342
rect 2625 -388 2779 -376
<< polycont >>
rect 571 -376 705 -342
rect 829 -376 963 -342
rect 1087 -376 1221 -342
rect 1345 -376 1479 -342
rect 1603 -376 1737 -342
rect 1861 -376 1995 -342
rect 2119 -376 2253 -342
rect 2377 -376 2511 -342
rect 2635 -376 2769 -342
<< locali >>
rect 190 1302 228 1324
rect 174 -12 244 1302
rect 2664 2 2734 1316
rect 2680 -12 2718 2
rect 22 -228 222 -206
rect -24 -236 10 -230
rect 22 -236 204 -228
rect -24 -376 206 -236
rect 2876 -238 3038 -204
rect 3072 -238 3106 -206
rect 561 -376 571 -342
rect 705 -376 715 -342
rect 819 -376 829 -342
rect 963 -376 973 -342
rect 1077 -376 1087 -342
rect 1221 -376 1231 -342
rect 1335 -376 1345 -342
rect 1479 -376 1489 -342
rect 1593 -376 1603 -342
rect 1737 -376 1747 -342
rect 1851 -376 1861 -342
rect 1995 -376 2005 -342
rect 2109 -376 2119 -342
rect 2253 -376 2263 -342
rect 2367 -376 2377 -342
rect 2511 -376 2521 -342
rect 2625 -376 2635 -342
rect 2769 -376 2779 -342
rect 2876 -376 3106 -238
rect -24 -448 10 -376
rect 3072 -436 3106 -376
rect -24 -1752 10 -1540
rect 3072 -1762 3106 -1550
<< viali >>
rect 380 1296 530 1332
rect 571 -376 705 -342
rect 829 -376 963 -342
rect 1087 -376 1221 -342
rect 1345 -376 1479 -342
rect 1603 -376 1737 -342
rect 1861 -376 1995 -342
rect 2119 -376 2253 -342
rect 2377 -376 2511 -342
rect 2635 -376 2769 -342
rect 1292 -1762 1670 -1728
<< metal1 >>
rect 350 1332 566 1410
rect 350 1296 380 1332
rect 530 1296 566 1332
rect 350 1290 566 1296
rect 350 1166 400 1290
rect 516 1166 566 1290
rect 682 1258 1230 1286
rect 682 1168 732 1258
rect 848 1202 1064 1230
rect 848 1166 898 1202
rect 1014 1166 1064 1202
rect 1180 1168 1230 1258
rect 1346 1260 1894 1288
rect 1346 1170 1396 1260
rect 1512 1202 1728 1230
rect 1512 1166 1562 1202
rect 1678 1166 1728 1202
rect 1844 1170 1894 1260
rect 2010 1258 2558 1286
rect 2010 1168 2060 1258
rect 2176 1202 2392 1230
rect 2176 1166 2226 1202
rect 2342 1166 2392 1202
rect 2508 1168 2558 1258
rect 350 50 400 130
rect 516 106 566 142
rect 682 132 686 134
rect 682 106 732 132
rect 516 78 732 106
rect 848 50 898 128
rect 350 22 898 50
rect 1014 52 1064 142
rect 1180 108 1230 144
rect 1346 108 1396 144
rect 1180 80 1396 108
rect 1512 52 1562 142
rect 1014 24 1562 52
rect 1678 50 1728 140
rect 1844 106 1894 142
rect 2010 106 2060 142
rect 1844 78 2060 106
rect 2176 50 2226 140
rect 1678 22 2226 50
rect 2342 -106 2392 158
rect 2508 -106 2558 164
rect 2342 -250 2558 -106
rect 234 -294 2850 -250
rect 234 -464 268 -294
rect 304 -332 456 -326
rect 304 -384 310 -332
rect 450 -384 456 -332
rect 562 -332 714 -326
rect 562 -336 568 -332
rect 561 -382 568 -336
rect 708 -336 714 -332
rect 304 -390 456 -384
rect 562 -384 568 -382
rect 708 -382 715 -336
rect 708 -384 714 -382
rect 562 -388 714 -384
rect 750 -462 784 -294
rect 820 -332 972 -326
rect 820 -336 826 -332
rect 819 -382 826 -336
rect 966 -336 972 -332
rect 1078 -332 1230 -326
rect 1078 -336 1084 -332
rect 820 -384 826 -382
rect 966 -382 973 -336
rect 1077 -382 1084 -336
rect 1224 -336 1230 -332
rect 966 -384 972 -382
rect 820 -388 972 -384
rect 1078 -384 1084 -382
rect 1224 -382 1231 -336
rect 1224 -384 1230 -382
rect 1078 -388 1230 -384
rect 1266 -462 1300 -294
rect 1336 -332 1488 -326
rect 1336 -336 1342 -332
rect 1335 -382 1342 -336
rect 1482 -336 1488 -332
rect 1594 -332 1746 -326
rect 1594 -336 1600 -332
rect 1336 -384 1342 -382
rect 1482 -382 1489 -336
rect 1593 -382 1600 -336
rect 1740 -336 1746 -332
rect 1482 -384 1488 -382
rect 1336 -388 1488 -384
rect 1594 -384 1600 -382
rect 1740 -382 1747 -336
rect 1740 -384 1746 -382
rect 1594 -388 1746 -384
rect 1782 -456 1816 -294
rect 1852 -332 2004 -326
rect 1852 -336 1858 -332
rect 1851 -382 1858 -336
rect 1998 -336 2004 -332
rect 2110 -332 2262 -326
rect 2110 -336 2116 -332
rect 1852 -384 1858 -382
rect 1998 -382 2005 -336
rect 2109 -382 2116 -336
rect 2256 -336 2262 -332
rect 1998 -384 2004 -382
rect 1852 -388 2004 -384
rect 2110 -384 2116 -382
rect 2256 -382 2263 -336
rect 2256 -384 2262 -382
rect 2110 -388 2262 -384
rect 2298 -456 2332 -294
rect 2368 -332 2520 -326
rect 2368 -336 2374 -332
rect 2367 -382 2374 -336
rect 2514 -336 2520 -332
rect 2626 -332 2778 -326
rect 2626 -336 2632 -332
rect 2368 -384 2374 -382
rect 2514 -382 2521 -336
rect 2625 -382 2632 -336
rect 2772 -336 2778 -332
rect 2514 -384 2520 -382
rect 2368 -388 2520 -384
rect 2626 -384 2632 -382
rect 2772 -382 2779 -336
rect 2772 -384 2778 -382
rect 2626 -388 2778 -384
rect 2816 -456 2850 -294
rect 492 -1710 526 -1502
rect 1008 -1710 1042 -1502
rect 1524 -1710 1558 -1514
rect 2040 -1710 2074 -1514
rect 2556 -1710 2590 -1506
rect 492 -1728 2590 -1710
rect 492 -1762 1292 -1728
rect 1670 -1762 2590 -1728
rect 492 -1772 2590 -1762
rect 1292 -1814 1670 -1772
<< via1 >>
rect 310 -384 450 -332
rect 568 -342 708 -332
rect 568 -376 571 -342
rect 571 -376 705 -342
rect 705 -376 708 -342
rect 568 -384 708 -376
rect 826 -342 966 -332
rect 826 -376 829 -342
rect 829 -376 963 -342
rect 963 -376 966 -342
rect 826 -384 966 -376
rect 1084 -342 1224 -332
rect 1084 -376 1087 -342
rect 1087 -376 1221 -342
rect 1221 -376 1224 -342
rect 1084 -384 1224 -376
rect 1342 -342 1482 -332
rect 1342 -376 1345 -342
rect 1345 -376 1479 -342
rect 1479 -376 1482 -342
rect 1342 -384 1482 -376
rect 1600 -342 1740 -332
rect 1600 -376 1603 -342
rect 1603 -376 1737 -342
rect 1737 -376 1740 -342
rect 1600 -384 1740 -376
rect 1858 -342 1998 -332
rect 1858 -376 1861 -342
rect 1861 -376 1995 -342
rect 1995 -376 1998 -342
rect 1858 -384 1998 -376
rect 2116 -342 2256 -332
rect 2116 -376 2119 -342
rect 2119 -376 2253 -342
rect 2253 -376 2256 -342
rect 2116 -384 2256 -376
rect 2374 -342 2514 -332
rect 2374 -376 2377 -342
rect 2377 -376 2511 -342
rect 2511 -376 2514 -342
rect 2374 -384 2514 -376
rect 2632 -342 2772 -332
rect 2632 -376 2635 -342
rect 2635 -376 2769 -342
rect 2769 -376 2772 -342
rect 2632 -384 2772 -376
<< metal2 >>
rect -360 -332 2778 -326
rect -360 -384 310 -332
rect 450 -384 568 -332
rect 708 -384 826 -332
rect 966 -384 1084 -332
rect 1224 -384 1342 -332
rect 1482 -384 1600 -332
rect 1740 -384 1858 -332
rect 1998 -384 2116 -332
rect 2256 -384 2374 -332
rect 2514 -384 2632 -332
rect 2772 -384 2778 -332
rect -360 -390 2778 -384
use sky130_fd_pr__nfet_g5v0d10v5_HLHUBB  sky130_fd_pr__nfet_g5v0d10v5_HLHUBB_0
timestamp 1693046372
transform 1 0 1541 0 1 -983
box -1747 -827 1747 827
use sky130_fd_pr__res_high_po_0p35_HS5UUT  sky130_fd_pr__res_high_po_0p35_HS5UUT_0
timestamp 1693010461
transform 1 0 1454 0 1 654
box -1507 -707 1507 707
<< labels >>
flabel metal1 350 1332 566 1410 0 FreeSans 320 0 0 0 VDD
port 1 nsew
flabel metal1 1292 -1814 1670 -1744 0 FreeSans 320 0 0 0 VSS
port 2 nsew
flabel metal2 -360 -390 310 -326 0 FreeSans 320 0 0 0 VIN
port 3 nsew
flabel metal1 2342 -294 2558 -106 0 FreeSans 320 0 0 0 VOUT
port 4 nsew
<< end >>
