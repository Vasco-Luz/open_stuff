magic
tech sky130A
magscale 1 2
timestamp 1693346665
<< locali >>
rect -456 4104 -416 4130
rect -472 3558 -400 4104
rect 2682 3558 2754 4104
rect -472 2828 -400 3360
rect -472 2820 -398 2828
rect -472 2812 312 2820
rect -456 2790 -416 2812
rect -400 1342 312 2812
rect 2682 2802 2756 3362
rect 2698 2794 2738 2802
rect -596 1114 -54 1188
rect 144 1114 698 1186
rect -608 782 -54 848
rect 144 782 698 854
<< viali >>
rect -290 4082 -90 4118
<< metal1 >>
rect -296 4118 -78 4150
rect -296 4082 -290 4118
rect -90 4082 -78 4118
rect -296 4074 -78 4082
rect -296 3564 -244 4074
rect -130 3564 -78 4074
rect 36 4066 586 4094
rect 36 3564 88 4066
rect 202 4008 420 4038
rect 202 3564 254 4008
rect 368 3564 420 4008
rect 534 3564 586 4066
rect 700 4066 1250 4094
rect 700 3564 752 4066
rect 866 4008 1084 4038
rect 866 3564 918 4008
rect 1032 3564 1084 4008
rect 1198 3564 1250 4066
rect 1364 4066 1914 4094
rect 1364 3564 1416 4066
rect 1530 4008 1748 4038
rect 1530 3564 1582 4008
rect 1696 3564 1748 4008
rect 1862 3564 1914 4066
rect 2028 4066 2578 4094
rect 2028 3564 2080 4066
rect 2194 4008 2412 4038
rect 2194 3564 2246 4008
rect 2360 3564 2412 4008
rect 2526 3564 2578 4066
rect -296 3058 -244 3354
rect -296 2946 -260 3058
rect -296 2852 -244 2946
rect -130 2910 -78 3354
rect 36 2910 90 3354
rect -130 2880 90 2910
rect 202 2852 254 3354
rect -296 2824 254 2852
rect 368 2852 422 3354
rect 534 2910 588 3354
rect 700 2910 754 3354
rect 534 2880 754 2910
rect 864 2852 918 3354
rect 368 2824 918 2852
rect 1032 2852 1086 3354
rect 1198 2910 1250 3354
rect 1364 2910 1416 3374
rect 1198 2880 1416 2910
rect 1530 2852 1584 3354
rect 1032 2824 1584 2852
rect 1696 2852 1750 3354
rect 1862 2910 1916 3354
rect 2028 2910 2082 3354
rect 1862 2880 2082 2910
rect 2192 2852 2246 3354
rect 1696 2824 2246 2852
rect 2360 2786 2414 3356
rect 2524 2786 2582 3354
rect 2360 2758 2582 2786
rect 2458 1742 2499 2758
rect 800 1010 866 1016
rect -734 958 -346 1010
rect 150 958 808 1010
rect 860 958 866 1010
rect 800 952 866 958
rect 2116 1010 2176 1016
rect 2116 952 2176 958
rect 2420 964 2430 1050
rect 2510 964 2520 1050
rect 2420 956 2520 964
<< via1 >>
rect 808 958 860 1010
rect 2116 958 2176 1010
rect 2430 964 2510 1050
<< metal2 >>
rect 800 1010 2184 1018
rect 800 958 808 1010
rect 860 958 2116 1010
rect 2176 958 2184 1010
rect 800 948 2184 958
rect 2420 964 2430 1050
rect 2510 964 2520 1050
rect 2420 956 2520 964
rect 2432 672 2508 956
rect 2432 -56 2510 672
use sky130_fd_pr__res_high_po_0p35_6HBKDU  sky130_fd_pr__res_high_po_0p35_6HBKDU_0
timestamp 1693271015
transform 1 0 1141 0 1 3459
box -1839 -707 1839 707
use sky130_fd_pr__res_high_po_0p35_8ZDV9T  sky130_fd_pr__res_high_po_0p35_8ZDV9T_0
timestamp 1693271449
transform 0 1 45 -1 0 984
box -428 -707 428 707
use sky130_fd_pr__rf_npn_05v5_W1p00L2p00  sky130_fd_pr__rf_npn_05v5_W1p00L2p00_0 ~/Desktop/pdk/sky130A/libs.ref/sky130_fd_pr/mag
timestamp 1692646696
transform 1 0 1594 0 1 6
box 0 0 1724 1924
<< labels >>
flabel metal1 -296 4118 -78 4150 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal2 2432 -56 2510 672 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 -734 958 -346 1010 0 FreeSans 1600 0 0 0 VIN
port 3 nsew
flabel metal1 2458 1742 2499 2786 0 FreeSans 1600 0 0 0 VOUT
port 4 nsew
<< end >>
